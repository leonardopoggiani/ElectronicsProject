library IEEE;
use IEEE.std_logic_1164.all;

entity fullAdder_tb is   
end fullAdder_tb;

architecture bhv of fullAdder_tb is 
   
	constant T_CLK   : time := 10 ns; 
	constant T_RESET : time := 25 ns; 
	
	signal a_tb		: std_logic := '0'; 
	signal b_tb		: std_logic := '0'; 
	signal c_i_tb	: std_logic := '0'; 
	signal o_tb		: std_logic; 		
	signal c_o_tb	: std_logic; 		
	
	signal clk_tb : std_logic := '0'; 
	signal rst_tb  : std_logic := '0'; 	
	signal end_sim : std_logic := '1';
  
    component fullAdder is   
		port(
                a   : in std_logic;
                b   : in std_logic;
                c_i : in std_logic;
                o   : out std_logic;
                c_o : out std_logic
	       );
	end component;
	
	
	begin
	
	  clk_tb <= (not(clk_tb) and end_sim) after T_CLK / 2;  
	  rst_tb <= '1' after T_RESET;
	  
	  test_fullAdder: fullAdder 
	   port map(
			a       => a_tb,
			b       => b_tb,
			c_i     => c_i_tb,
	        o 	=> o_tb,
			c_o		=> c_o_tb
		);
	  

	  
	  d_process: process(clk_tb, rst_tb) 
		variable t : integer := 0;
	  begin
	    if(rst_tb = '0') then
		  a_tb 	<= '0';
		  b_tb 	<= '0';
		  c_i_tb 	<= '0';	
		  t := 0;
		elsif(rising_edge(clk_tb)) then
		  case(t) is  
		    when 1 => a_tb <= '0'; b_tb <= '0';
			
			when 2 => a_tb <= '0'; b_tb <= '1';
			
			when 3 => a_tb <= '1'; b_tb <= '0';
			
			when 4 => a_tb <= '1'; b_tb <= '1';
			
			when 10 => end_sim <= '0'; 
            when others => null;
			
		  end case;
		  t := t + 1; 
		end if;
	  end process;
	
end bhv;
