library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all; -- for the casting 
	
-- This testbench aims to check if the output
-- of the filter is the same as the one designed in MATLAB

entity IIR_TB_Synth is
end IIR_TB_Synth;

architecture TB_Arch of IIR_TB_Synth is	

component IIR  
	generic (Nbit : natural := 8);
	port (
		clk		:	in	std_logic;
		rst_l	:	in	std_logic;
		x		:	in	std_logic_vector(Nbit-1 downto 0);	
		y		:	out	std_logic_vector(Nbit-1 downto 0)
	);
end component;

	constant BITS		:	natural	:=	16;
	constant SAMPLES 	:	natural	:= 	1000;

	signal clk		: 	std_logic	:= '0'; 
	signal rst_l 	: 	std_logic;
	signal sample	:	std_logic_vector(BITS-1 downto 0);
	signal output	:	std_logic_vector(BITS-1 downto 0);
	signal expected	:	std_logic_vector(BITS-1 downto 0);
	
	signal enable	:	std_logic	:=	'1';
	
	-- Data type to store the sequence of samples
	type WAV_IN is array (0 to SAMPLES-1) of std_logic_vector(BITS-1 downto 0);

begin
	
	filter: IIR
	generic map(BITS)
	port map(clk, rst_l, sample, output);
	
	-- clock generator
	clk <= not clk and enable after 11338 ns; -- 44100Hz clock
	
	-- stimuli
	driver_p: process
	
	variable input : WAV_IN := ("0000000000000000",
								"0000000000000000",
								"1111111111111111",
								"1111111111111110",
								"1111111111111111",
								"1111111111111111",
								"1111111111111110",
								"0000000000000000",
								"0000000000000010",
								"0000000000000000",
								"1111111111111111",
								"0000000000000000",
								"0000000000000000",
								"1111111111111111",
								"1111111111111110",
								"0000000000000000",
								"1111111111111111",
								"1111111111111110",
								"1111111111111110",
								"1111111111111111",
								"1111111111111110",
								"1111111111111111",
								"0000000000000000",
								"1111111111111111",
								"1111111111111111",
								"0000000000000000",
								"1111111111111111",
								"1111111111111110",
								"1111111111111111",
								"1111111111111111",
								"1111111111111111",
								"0000000000000000",
								"1111111111111110",
								"1111111111111111",
								"0000000000000000",
								"0000000000000001",
								"0000000000000000",
								"0000000000000000",
								"1111111111111111",
								"0000000000000000",
								"1111111111111111",
								"1111111111111111",
								"0000000000000000",
								"0000000000000000",
								"1111111111111111",
								"1111111111111111",
								"0000000000000000",
								"0000000000000001",
								"0000000000000001",
								"0000000000000001",
								"0000000000000000",
								"0000000000000000",
								"0000000000000001",
								"1111111111111111",
								"1111111111111110",
								"0000000000000000",
								"0000000000000000",
								"1111111111111111",
								"0000000000000000",
								"1111111111111111",
								"1111111111111111",
								"0000000000000000",
								"1111111111111111",
								"1111111111111111",
								"0000000000000000",
								"1111111111111111",
								"1111111111111111",
								"0000000000000000",
								"0000000000000000",
								"1111111111111111",
								"1111111111111111",
								"1111111111111110",
								"1111111111111111",
								"1111111111111111",
								"1111111111111110",
								"1111111111111111",
								"0000000000000000",
								"1111111111111111",
								"1111111111111111",
								"1111111111111111",
								"1111111111111111",
								"0000000000000001",
								"0000000000000010",
								"0000000000000000",
								"1111111111111111",
								"1111111111111111",
								"1111111111111111",
								"1111111111111111",
								"1111111111111111",
								"0000000000000000",
								"0000000000000000",
								"1111111111111111",
								"1111111111111111",
								"0000000000000000",
								"1111111111111111",
								"1111111111111110",
								"1111111111111111",
								"1111111111111111",
								"0000000000000000",
								"0000000000000000",
								"0000000000000000",
								"0000000000000000",
								"1111111111111110",
								"1111111111111111",
								"1111111111111111",
								"0000000000000000",
								"1111111111111111",
								"0000000000000001",
								"0000000000000000",
								"1111111111111111",
								"0000000000000000",
								"0000000000000001",
								"1111111111111111",
								"0000000000000000",
								"0000000000000001",
								"0000000000000001",
								"0000000000000000",
								"0000000000000000",
								"0000000000000000",
								"0000000000000000",
								"1111111111111111",
								"1111111111111111",
								"0000000000000000",
								"0000000000000000",
								"0000000000000000",
								"0000000000000000",
								"1111111111111111",
								"1111111111111111",
								"1111111111111111",
								"0000000000000000",
								"1111111111111111",
								"0000000000000000",
								"1111111111111110",
								"1111111111111110",
								"0000000000000000",
								"0000000000000000",
								"1111111111111110",
								"1111111111111101",
								"1111111111111111",
								"1111111111111111",
								"1111111111111111",
								"1111111111111110",
								"1111111111111111",
								"0000000000000000",
								"1111111111111111",
								"1111111111111111",
								"1111111111111110",
								"1111111111111111",
								"0000000000000001",
								"0000000000000000",
								"1111111111111111",
								"1111111111111111",
								"0000000000000000",
								"1111111111111111",
								"1111111111111111",
								"1111111111111111",
								"1111111111111111",
								"1111111111111111",
								"0000000000000000",
								"1111111111111111",
								"1111111111111101",
								"1111111111111110",
								"1111111111111111",
								"0000000000000000",
								"0000000000000000",
								"1111111111111111",
								"1111111111111111",
								"1111111111111111",
								"1111111111111110",
								"1111111111111111",
								"0000000000000000",
								"0000000000000000",
								"1111111111111111",
								"1111111111111110",
								"1111111111111110",
								"1111111111111111",
								"0000000000000000",
								"0000000000000000",
								"0000000000000000",
								"1111111111111111",
								"1111111111111111",
								"0000000000000000",
								"0000000000000000",
								"1111111111111111",
								"1111111111111111",
								"0000000000000000",
								"0000000000000000",
								"1111111111111111",
								"0000000000000000",
								"1111111111111111",
								"1111111111111110",
								"1111111111111101",
								"1111111111111111",
								"1111111111111111",
								"1111111111111111",
								"0000000000000001",
								"0000000000000000",
								"0000000000000000",
								"0000000000000000",
								"0000000000000000",
								"1111111111111111",
								"1111111111111111",
								"1111111111111111",
								"1111111111111111",
								"1111111111111110",
								"1111111111111110",
								"0000000000000000",
								"0000000000000000",
								"1111111111111110",
								"1111111111111111",
								"0000000000000001",
								"0000000000000000",
								"1111111111111101",
								"1111111111111110",
								"1111111111111110",
								"1111111111111110",
								"1111111111111111",
								"1111111111111111",
								"1111111111111110",
								"1111111111111110",
								"1111111111111110",
								"1111111111111110",
								"1111111111111110",
								"1111111111111101",
								"1111111111111111",
								"1111111111111111",
								"1111111111111111",
								"0000000000000000",
								"1111111111111111",
								"1111111111111110",
								"1111111111111111",
								"0000000000000000",
								"1111111111111111",
								"1111111111111111",
								"1111111111111111",
								"1111111111111111",
								"1111111111111111",
								"0000000000000000",
								"0000000000000000",
								"0000000000000000",
								"1111111111111111",
								"1111111111111110",
								"1111111111111111",
								"0000000000000000",
								"1111111111111111",
								"0000000000000000",
								"0000000000000000",
								"1111111111111111",
								"1111111111111111",
								"1111111111111110",
								"1111111111111110",
								"1111111111111111",
								"1111111111111110",
								"1111111111111111",
								"0000000000000001",
								"0000000000000000",
								"1111111111111111",
								"1111111111111111",
								"1111111111111111",
								"1111111111111111",
								"1111111111111111",
								"1111111111111111",
								"1111111111111111",
								"0000000000000000",
								"0000000000000010",
								"0000000000000001",
								"0000000000000000",
								"1111111111111110",
								"1111111111111111",
								"0000000000000000",
								"0000000000000000",
								"0000000000000000",
								"0000000000000000",
								"1111111111111111",
								"1111111111111111",
								"1111111111111110",
								"1111111111111101",
								"1111111111111110",
								"1111111111111110",
								"1111111111111110",
								"1111111111111110",
								"0000000000000000",
								"1111111111111111",
								"1111111111111111",
								"1111111111111110",
								"1111111111111110",
								"1111111111111111",
								"1111111111111111",
								"1111111111111111",
								"1111111111111111",
								"1111111111111111",
								"1111111111111110",
								"1111111111111101",
								"1111111111111111",
								"1111111111111111",
								"1111111111111111",
								"1111111111111110",
								"1111111111111111",
								"0000000000000000",
								"1111111111111110",
								"1111111111111110",
								"1111111111111111",
								"1111111111111111",
								"1111111111111110",
								"0000000000000000",
								"0000000000000000",
								"1111111111111111",
								"0000000000000000",
								"0000000000000000",
								"1111111111111111",
								"1111111111111110",
								"1111111111111111",
								"0000000000000000",
								"1111111111111111",
								"1111111111111111",
								"1111111111111101",
								"1111111111111101",
								"1111111111111110",
								"1111111111111111",
								"1111111111111110",
								"1111111111111111",
								"1111111111111111",
								"0000000000000000",
								"0000000000000000",
								"1111111111111111",
								"1111111111111111",
								"1111111111111111",
								"0000000000000000",
								"1111111111111111",
								"1111111111111111",
								"1111111111111111",
								"0000000000000000",
								"1111111111111111",
								"0000000000000000",
								"1111111111111111",
								"1111111111111111",
								"1111111111111111",
								"1111111111111111",
								"1111111111111111",
								"1111111111111110",
								"1111111111111111",
								"0000000000000001",
								"0000000000000000",
								"1111111111111110",
								"0000000000000000",
								"0000000000000000",
								"1111111111111111",
								"1111111111111111",
								"1111111111111111",
								"1111111111111101",
								"1111111111111110",
								"1111111111111111",
								"1111111111111111",
								"1111111111111111",
								"0000000000000001",
								"0000000000000010",
								"0000000000000000",
								"1111111111111111",
								"1111111111111111",
								"0000000000000000",
								"1111111111111110",
								"1111111111111110",
								"0000000000000000",
								"1111111111111111",
								"1111111111111110",
								"0000000000000000",
								"1111111111111111",
								"1111111111111111",
								"0000000000000000",
								"1111111111111111",
								"1111111111111110",
								"1111111111111111",
								"0000000000000000",
								"1111111111111111",
								"0000000000000000",
								"0000000000000000",
								"1111111111111111",
								"1111111111111110",
								"1111111111111111",
								"0000000000000001",
								"0000000000000001",
								"0000000000000001",
								"0000000000000000",
								"0000000000000001",
								"0000000000000001",
								"0000000000000001",
								"0000000000000000",
								"1111111111111111",
								"0000000000000001",
								"0000000000000000",
								"1111111111111111",
								"1111111111111111",
								"1111111111111111",
								"1111111111111111",
								"1111111111111110",
								"1111111111111110",
								"1111111111111111",
								"1111111111111111",
								"1111111111111111",
								"1111111111111111",
								"1111111111111111",
								"1111111111111111",
								"0000000000000000",
								"1111111111111111",
								"1111111111111110",
								"1111111111111111",
								"1111111111111111",
								"1111111111111110",
								"1111111111111110",
								"0000000000000000",
								"0000000000000000",
								"1111111111111111",
								"1111111111111111",
								"1111111111111111",
								"1111111111111111",
								"1111111111111111",
								"1111111111111110",
								"1111111111111110",
								"1111111111111111",
								"1111111111111110",
								"1111111111111110",
								"1111111111111111",
								"0000000000000000",
								"0000000000000000",
								"0000000000000000",
								"1111111111111111",
								"1111111111111111",
								"0000000000000000",
								"1111111111111111",
								"1111111111111111",
								"1111111111111110",
								"1111111111111101",
								"1111111111111101",
								"1111111111111101",
								"1111111111111101",
								"1111111111111110",
								"1111111111111110",
								"1111111111111110",
								"1111111111111110",
								"1111111111111111",
								"0000000000000000",
								"1111111111111111",
								"1111111111111111",
								"1111111111111111",
								"0000000000000000",
								"0000000000000001",
								"0000000000000000",
								"1111111111111111",
								"1111111111111110",
								"1111111111111110",
								"0000000000000000",
								"1111111111111111",
								"0000000000000000",
								"0000000000000000",
								"1111111111111111",
								"1111111111111110",
								"0000000000000000",
								"0000000000000001",
								"1111111111111111",
								"0000000000000000",
								"0000000000000000",
								"0000000000000000",
								"0000000000000000",
								"1111111111111111",
								"1111111111111111",
								"0000000000000000",
								"0000000000000000",
								"1111111111111111",
								"0000000000000000",
								"1111111111111111",
								"1111111111111111",
								"1111111111111111",
								"1111111111111111",
								"1111111111111111",
								"0000000000000000",
								"1111111111111111",
								"1111111111111111",
								"0000000000000000",
								"0000000000000000",
								"1111111111111111",
								"0000000000000000",
								"0000000000000001",
								"1111111111111111",
								"0000000000000000",
								"0000000000000000",
								"1111111111111111",
								"1111111111111111",
								"0000000000000000",
								"0000000000000000",
								"0000000000000001",
								"0000000000000001",
								"0000000000000000",
								"1111111111111111",
								"1111111111111111",
								"1111111111111111",
								"0000000000000000",
								"1111111111111111",
								"1111111111111110",
								"1111111111111111",
								"1111111111111111",
								"1111111111111111",
								"0000000000000001",
								"0000000000000001",
								"1111111111111111",
								"1111111111111111",
								"0000000000000000",
								"0000000000000000",
								"0000000000000000",
								"1111111111111111",
								"1111111111111111",
								"0000000000000001",
								"0000000000000000",
								"1111111111111111",
								"1111111111111110",
								"0000000000000000",
								"1111111111111111",
								"1111111111111111",
								"0000000000000000",
								"1111111111111111",
								"1111111111111111",
								"0000000000000001",
								"1111111111111111",
								"1111111111111111",
								"1111111111111111",
								"1111111111111111",
								"0000000000000000",
								"0000000000000001",
								"1111111111111111",
								"0000000000000000",
								"0000000000000000",
								"1111111111111111",
								"1111111111111111",
								"0000000000000000",
								"0000000000000000",
								"0000000000000000",
								"1111111111111111",
								"1111111111111111",
								"0000000000000001",
								"0000000000000000",
								"1111111111111111",
								"1111111111111111",
								"1111111111111110",
								"1111111111111101",
								"1111111111111111",
								"0000000000000000",
								"1111111111111110",
								"1111111111111110",
								"1111111111111111",
								"1111111111111111",
								"1111111111111110",
								"1111111111111110",
								"1111111111111110",
								"1111111111111111",
								"1111111111111111",
								"1111111111111110",
								"1111111111111110",
								"1111111111111110",
								"1111111111111111",
								"1111111111111111",
								"1111111111111111",
								"1111111111111110",
								"0000000000000000",
								"1111111111111111",
								"1111111111111111",
								"0000000000000000",
								"0000000000000000",
								"0000000000000000",
								"0000000000000000",
								"1111111111111111",
								"0000000000000000",
								"1111111111111111",
								"1111111111111111",
								"0000000000000001",
								"0000000000000000",
								"1111111111111111",
								"1111111111111111",
								"0000000000000000",
								"1111111111111111",
								"1111111111111110",
								"1111111111111110",
								"1111111111111111",
								"1111111111111111",
								"1111111111111111",
								"1111111111111111",
								"0000000000000000",
								"1111111111111111",
								"1111111111111110",
								"1111111111111110",
								"1111111111111110",
								"1111111111111110",
								"1111111111111110",
								"1111111111111111",
								"0000000000000001",
								"0000000000000001",
								"0000000000000000",
								"1111111111111111",
								"1111111111111111",
								"1111111111111110",
								"1111111111111110",
								"1111111111111111",
								"0000000000000000",
								"1111111111111111",
								"1111111111111110",
								"1111111111111111",
								"1111111111111111",
								"1111111111111111",
								"0000000000000000",
								"0000000000000001",
								"0000000000000000",
								"1111111111111101",
								"1111111111111111",
								"0000000000000000",
								"1111111111111110",
								"1111111111111111",
								"0000000000000000",
								"1111111111111111",
								"1111111111111111",
								"0000000000000000",
								"0000000000000000",
								"1111111111111111",
								"1111111111111111",
								"1111111111111111",
								"1111111111111111",
								"1111111111111110",
								"1111111111111110",
								"0000000000000000",
								"1111111111111111",
								"1111111111111101",
								"1111111111111110",
								"1111111111111111",
								"1111111111111101",
								"0000000000000000",
								"0000000000000000",
								"1111111111111111",
								"1111111111111111",
								"0000000000000000",
								"1111111111111111",
								"1111111111111111",
								"1111111111111111",
								"1111111111111111",
								"1111111111111111",
								"1111111111111111",
								"0000000000000000",
								"1111111111111111",
								"0000000000000000",
								"1111111111111111",
								"1111111111111111",
								"1111111111111111",
								"1111111111111111",
								"1111111111111111",
								"1111111111111111",
								"0000000000000000",
								"0000000000000001",
								"0000000000000000",
								"1111111111111111",
								"1111111111111111",
								"1111111111111111",
								"1111111111111111",
								"0000000000000000",
								"0000000000000000",
								"0000000000000000",
								"0000000000000000",
								"1111111111111111",
								"0000000000000000",
								"0000000000000001",
								"0000000000000000",
								"0000000000000000",
								"0000000000000001",
								"0000000000000000",
								"1111111111111111",
								"1111111111111111",
								"1111111111111111",
								"0000000000000001",
								"0000000000000000",
								"1111111111111111",
								"1111111111111111",
								"1111111111111111",
								"0000000000000000",
								"0000000000000000",
								"1111111111111111",
								"0000000000000000",
								"0000000000000000",
								"1111111111111111",
								"1111111111111111",
								"1111111111111110",
								"1111111111111111",
								"0000000000000000",
								"0000000000000000",
								"1111111111111110",
								"1111111111111110",
								"1111111111111111",
								"1111111111111111",
								"1111111111111111",
								"1111111111111111",
								"0000000000000000",
								"1111111111111111",
								"1111111111111110",
								"1111111111111110",
								"0000000000000000",
								"1111111111111111",
								"1111111111111101",
								"1111111111111111",
								"0000000000000000",
								"1111111111111110",
								"1111111111111111",
								"1111111111111111",
								"1111111111111110",
								"0000000000000000",
								"0000000000000001",
								"1111111111111111",
								"1111111111111111",
								"1111111111111111",
								"1111111111111110",
								"1111111111111111",
								"0000000000000000",
								"1111111111111111",
								"1111111111111111",
								"1111111111111111",
								"1111111111111111",
								"0000000000000000",
								"0000000000000000",
								"1111111111111111",
								"0000000000000001",
								"0000000000000001",
								"1111111111111110",
								"1111111111111111",
								"0000000000000000",
								"1111111111111110",
								"1111111111111101",
								"1111111111111110",
								"0000000000000000",
								"1111111111111110",
								"1111111111111110",
								"1111111111111111",
								"1111111111111111",
								"1111111111111111",
								"1111111111111111",
								"1111111111111111",
								"1111111111111111",
								"0000000000000000",
								"0000000000000000",
								"1111111111111111",
								"1111111111111111",
								"1111111111111111",
								"0000000000000000",
								"0000000000000000",
								"1111111111111111",
								"0000000000000000",
								"0000000000000000",
								"0000000000000000",
								"0000000000000000",
								"1111111111111111",
								"1111111111111110",
								"1111111111111101",
								"0000000000000000",
								"0000000000000000",
								"1111111111111110",
								"0000000000000000",
								"0000000000000000",
								"0000000000000000",
								"0000000000000000",
								"0000000000000000",
								"1111111111111111",
								"0000000000000000",
								"0000000000000000",
								"1111111111111111",
								"1111111111111111",
								"1111111111111110",
								"1111111111111110",
								"1111111111111111",
								"1111111111111111",
								"1111111111111111",
								"0000000000000000",
								"1111111111111111",
								"1111111111111101",
								"1111111111111110",
								"1111111111111111",
								"1111111111111111",
								"1111111111111111",
								"0000000000000000",
								"1111111111111111",
								"0000000000000000",
								"0000000000000000",
								"1111111111111111",
								"0000000000000000",
								"0000000000000000",
								"1111111111111111",
								"1111111111111111",
								"0000000000000000",
								"0000000000000000",
								"0000000000000000",
								"0000000000000000",
								"0000000000000000",
								"0000000000000000",
								"1111111111111111",
								"1111111111111111",
								"0000000000000000",
								"1111111111111111",
								"1111111111111110",
								"1111111111111111",
								"0000000000000000",
								"1111111111111110",
								"1111111111111110",
								"1111111111111111",
								"1111111111111111",
								"1111111111111111",
								"1111111111111111",
								"1111111111111111",
								"1111111111111111",
								"1111111111111110",
								"1111111111111110",
								"1111111111111111",
								"1111111111111111",
								"0000000000000000",
								"1111111111111111",
								"1111111111111111",
								"0000000000000000",
								"0000000000000001",
								"0000000000000000",
								"1111111111111111",
								"0000000000000000",
								"1111111111111111",
								"1111111111111111",
								"1111111111111111",
								"1111111111111110",
								"1111111111111111",
								"1111111111111111",
								"0000000000000000",
								"0000000000000001",
								"0000000000000000",
								"0000000000000000",
								"0000000000000000",
								"1111111111111111",
								"0000000000000001",
								"0000000000000000",
								"1111111111111111",
								"1111111111111111",
								"0000000000000000",
								"0000000000000000",
								"0000000000000000",
								"1111111111111111",
								"1111111111111111",
								"1111111111111110",
								"1111111111111110",
								"1111111111111111",
								"0000000000000000",
								"0000000000000000",
								"1111111111111110",
								"1111111111111111",
								"1111111111111110",
								"1111111111111111",
								"0000000000000000",
								"0000000000000000",
								"1111111111111111",
								"0000000000000000",
								"1111111111111111",
								"1111111111111111",
								"1111111111111111",
								"0000000000000000",
								"1111111111111111",
								"1111111111111111",
								"1111111111111111",
								"0000000000000000",
								"0000000000000000",
								"0000000000000000",
								"1111111111111111",
								"1111111111111110",
								"1111111111111111",
								"1111111111111110",
								"1111111111111111",
								"1111111111111110",
								"1111111111111111",
								"1111111111111110",
								"1111111111111110",
								"1111111111111111",
								"1111111111111110",
								"1111111111111101",
								"1111111111111111",
								"1111111111111111",
								"1111111111111110",
								"0000000000000000",
								"0000000000000000",
								"1111111111111110",
								"1111111111111110",
								"1111111111111111",
								"1111111111111110",
								"1111111111111110",
								"1111111111111111",
								"1111111111111111",
								"1111111111111110",
								"1111111111111111",
								"1111111111111111",
								"1111111111111101",
								"1111111111111110",
								"1111111111111111",
								"1111111111111111",
								"1111111111111111",
								"0000000000000000",
								"0000000000000000",
								"1111111111111111",
								"1111111111111110",
								"1111111111111110",
								"0000000000000000",
								"0000000000000001",
								"0000000000000000",
								"1111111111111111",
								"1111111111111110",
								"1111111111111101",
								"0000000000000000",
								"0000000000000000",
								"1111111111111110",
								"1111111111111110",
								"1111111111111110",
								"1111111111111111",
								"0000000000000001",
								"0000000000000001",
								"1111111111111111",
								"1111111111111110",
								"1111111111111111",
								"1111111111111111",
								"1111111111111111",
								"0000000000000000",
								"1111111111111111",
								"1111111111111111",
								"0000000000000001",
								"0000000000000000",
								"1111111111111111",
								"0000000000000000",
								"0000000000000001",
								"1111111111111111",
								"1111111111111111",
								"0000000000000000",
								"0000000000000001",
								"0000000000000001",
								"1111111111111111",
								"1111111111111110",
								"0000000000000000",
								"0000000000000000",
								"1111111111111110",
								"0000000000000000",
								"0000000000000000",
								"1111111111111110",
								"1111111111111111",
								"0000000000000000",
								"1111111111111111",
								"1111111111111111",
								"1111111111111101",
								"1111111111111110",
								"1111111111111111",
								"0000000000000000",
								"1111111111111111",
								"1111111111111111",
								"0000000000000000",
								"0000000000000000",
								"0000000000000000",
								"1111111111111111",
								"1111111111111110",
								"1111111111111110",
								"0000000000000000",
								"0000000000000000",
								"1111111111111111",
								"0000000000000000",
								"0000000000000000",
								"1111111111111111",
								"0000000000000000",
								"0000000000000000",
								"1111111111111110",
								"0000000000000000",
								"0000000000000001",
								"0000000000000000",
								"1111111111111111",
								"1111111111111111",
								"1111111111111111",
								"0000000000000000",
								"0000000000000000",
								"1111111111111111",
								"1111111111111111",
								"0000000000000000",
								"1111111111111111",
								"1111111111111110",
								"1111111111111111",
								"1111111111111110",
								"1111111111111111",
								"0000000000000001",
								"0000000000000000",
								"1111111111111111",
								"1111111111111111",
								"1111111111111110",
								"1111111111111111",
								"0000000000000000",
								"1111111111111111",
								"1111111111111111",
								"1111111111111111",
								"1111111111111111",
								"0000000000000000",
								"1111111111111111",
								"1111111111111111",
								"0000000000000000",
								"0000000000000001",
								"1111111111111110"
								);
								
	variable expected_out : WAV_IN := ("0000000000000000",
										"0000000000000000",
										"0000000000000001",
										"0000000000000011",
										"0000000000000100",
										"0000000000000101",
										"0000000000000110",
										"0000000000000100",
										"0000000000000001",
										"0000000000000000",
										"1111111111111111",
										"1111111111111111",
										"0000000000000001",
										"0000000000000010",
										"0000000000000011",
										"0000000000000011",
										"0000000000000100",
										"0000000000000101",
										"0000000000000101",
										"0000000000000110",
										"0000000000000111",
										"0000000000000110",
										"0000000000000100",
										"0000000000000100",
										"0000000000000011",
										"0000000000000010",
										"0000000000000011",
										"0000000000000100",
										"0000000000000100",
										"0000000000000101",
										"0000000000000101",
										"0000000000000011",
										"0000000000000100",
										"0000000000000100",
										"0000000000000011",
										"0000000000000010",
										"0000000000000000",
										"1111111111111111",
										"0000000000000000",
										"0000000000000001",
										"0000000000000010",
										"0000000000000011",
										"0000000000000010",
										"0000000000000010",
										"0000000000000010",
										"0000000000000010",
										"0000000000000010",
										"0000000000000001",
										"1111111111111111",
										"1111111111111101",
										"1111111111111101",
										"1111111111111110",
										"1111111111111110",
										"0000000000000000",
										"0000000000000010",
										"0000000000000010",
										"0000000000000011",
										"0000000000000011",
										"0000000000000001",
										"0000000000000010",
										"0000000000000011",
										"0000000000000010",
										"0000000000000011",
										"0000000000000011",
										"0000000000000010",
										"0000000000000011",
										"0000000000000011",
										"0000000000000010",
										"0000000000000010",
										"0000000000000010",
										"0000000000000010",
										"0000000000000100",
										"0000000000000101",
										"0000000000000101",
										"0000000000000110",
										"0000000000000101",
										"0000000000000100",
										"0000000000000100",
										"0000000000000011",
										"0000000000000011",
										"0000000000000100",
										"0000000000000010",
										"1111111111111111",
										"1111111111111110",
										"1111111111111110",
										"0000000000000000",
										"0000000000000011",
										"0000000000000100",
										"0000000000000100",
										"0000000000000011",
										"0000000000000010",
										"0000000000000010",
										"0000000000000010",
										"0000000000000010",
										"0000000000000011",
										"0000000000000100",
										"0000000000000100",
										"0000000000000101",
										"0000000000000100",
										"0000000000000010",
										"0000000000000001",
										"0000000000000000",
										"0000000000000010",
										"0000000000000011",
										"0000000000000100",
										"0000000000000100",
										"0000000000000011",
										"0000000000000001",
										"0000000000000000",
										"0000000000000001",
										"0000000000000000",
										"0000000000000000",
										"0000000000000001",
										"0000000000000000",
										"1111111111111111",
										"1111111111111111",
										"1111111111111110",
										"1111111111111110",
										"1111111111111111",
										"0000000000000000",
										"0000000000000001",
										"0000000000000010",
										"0000000000000010",
										"0000000000000010",
										"0000000000000001",
										"0000000000000000",
										"0000000000000001",
										"0000000000000010",
										"0000000000000011",
										"0000000000000011",
										"0000000000000011",
										"0000000000000010",
										"0000000000000011",
										"0000000000000101",
										"0000000000000100",
										"0000000000000100",
										"0000000000000100",
										"0000000000000101",
										"0000000000000110",
										"0000000000000111",
										"0000000000000110",
										"0000000000000101",
										"0000000000000101",
										"0000000000000100",
										"0000000000000100",
										"0000000000000011",
										"0000000000000100",
										"0000000000000101",
										"0000000000000011",
										"0000000000000010",
										"0000000000000001",
										"0000000000000001",
										"0000000000000010",
										"0000000000000011",
										"0000000000000011",
										"0000000000000011",
										"0000000000000100",
										"0000000000000100",
										"0000000000000011",
										"0000000000000011",
										"0000000000000101",
										"0000000000000110",
										"0000000000000111",
										"0000000000000110",
										"0000000000000011",
										"0000000000000010",
										"0000000000000010",
										"0000000000000011",
										"0000000000000101",
										"0000000000000101",
										"0000000000000100",
										"0000000000000011",
										"0000000000000010",
										"0000000000000011",
										"0000000000000101",
										"0000000000000110",
										"0000000000000101",
										"0000000000000011",
										"0000000000000001",
										"0000000000000001",
										"0000000000000010",
										"0000000000000010",
										"0000000000000010",
										"0000000000000010",
										"0000000000000010",
										"0000000000000010",
										"0000000000000010",
										"0000000000000010",
										"0000000000000001",
										"0000000000000010",
										"0000000000000100",
										"0000000000000110",
										"0000000000000111",
										"0000000000000111",
										"0000000000000110",
										"0000000000000010",
										"0000000000000001",
										"0000000000000000",
										"1111111111111111",
										"0000000000000000",
										"0000000000000001",
										"0000000000000010",
										"0000000000000011",
										"0000000000000100",
										"0000000000000101",
										"0000000000000110",
										"0000000000000101",
										"0000000000000100",
										"0000000000000100",
										"0000000000000011",
										"0000000000000010",
										"0000000000000010",
										"0000000000000011",
										"0000000000000100",
										"0000000000000111",
										"0000000000001001",
										"0000000000000111",
										"0000000000000110",
										"0000000000000110",
										"0000000000000110",
										"0000000000000111",
										"0000000000001000",
										"0000000000001000",
										"0000000000001001",
										"0000000000001000",
										"0000000000000111",
										"0000000000000110",
										"0000000000000011",
										"0000000000000011",
										"0000000000000100",
										"0000000000000100",
										"0000000000000100",
										"0000000000000100",
										"0000000000000011",
										"0000000000000011",
										"0000000000000100",
										"0000000000000100",
										"0000000000000011",
										"0000000000000010",
										"0000000000000001",
										"0000000000000001",
										"0000000000000011",
										"0000000000000100",
										"0000000000000100",
										"0000000000000100",
										"0000000000000010",
										"0000000000000001",
										"0000000000000010",
										"0000000000000010",
										"0000000000000100",
										"0000000000000110",
										"0000000000000110",
										"0000000000000111",
										"0000000000000110",
										"0000000000000011",
										"0000000000000010",
										"0000000000000001",
										"0000000000000001",
										"0000000000000011",
										"0000000000000100",
										"0000000000000100",
										"0000000000000100",
										"0000000000000100",
										"0000000000000011",
										"0000000000000000",
										"1111111111111110",
										"1111111111111101",
										"1111111111111111",
										"0000000000000010",
										"0000000000000011",
										"0000000000000011",
										"0000000000000001",
										"0000000000000000",
										"0000000000000001",
										"0000000000000010",
										"0000000000000100",
										"0000000000000111",
										"0000000000001000",
										"0000000000001001",
										"0000000000001001",
										"0000000000001000",
										"0000000000000110",
										"0000000000000101",
										"0000000000000100",
										"0000000000000100",
										"0000000000000110",
										"0000000000000110",
										"0000000000000110",
										"0000000000000101",
										"0000000000000100",
										"0000000000000100",
										"0000000000000101",
										"0000000000000111",
										"0000000000000111",
										"0000000000000111",
										"0000000000000110",
										"0000000000000101",
										"0000000000000101",
										"0000000000000100",
										"0000000000000101",
										"0000000000000101",
										"0000000000000101",
										"0000000000000110",
										"0000000000000110",
										"0000000000000100",
										"0000000000000011",
										"0000000000000011",
										"0000000000000001",
										"0000000000000001",
										"0000000000000010",
										"0000000000000011",
										"0000000000000100",
										"0000000000000100",
										"0000000000000100",
										"0000000000000011",
										"0000000000000101",
										"0000000000001000",
										"0000000000001001",
										"0000000000001001",
										"0000000000001000",
										"0000000000000110",
										"0000000000000101",
										"0000000000000100",
										"0000000000000010",
										"0000000000000010",
										"0000000000000010",
										"0000000000000011",
										"0000000000000011",
										"0000000000000011",
										"0000000000000011",
										"0000000000000011",
										"0000000000000011",
										"0000000000000011",
										"0000000000000010",
										"0000000000000010",
										"0000000000000011",
										"0000000000000011",
										"0000000000000100",
										"0000000000000100",
										"0000000000000101",
										"0000000000000101",
										"0000000000000011",
										"0000000000000010",
										"0000000000000010",
										"0000000000000001",
										"0000000000000010",
										"0000000000000011",
										"0000000000000010",
										"0000000000000011",
										"0000000000000110",
										"0000000000000111",
										"0000000000000111",
										"0000000000000111",
										"0000000000000101",
										"0000000000000010",
										"1111111111111111",
										"1111111111111110",
										"1111111111111110",
										"0000000000000000",
										"0000000000000010",
										"0000000000000100",
										"0000000000000101",
										"0000000000000100",
										"0000000000000101",
										"0000000000000101",
										"0000000000000011",
										"0000000000000100",
										"0000000000000100",
										"0000000000000010",
										"0000000000000011",
										"0000000000000100",
										"0000000000000100",
										"0000000000000100",
										"0000000000000100",
										"0000000000000010",
										"0000000000000001",
										"0000000000000010",
										"0000000000000011",
										"0000000000000100",
										"0000000000000011",
										"0000000000000001",
										"1111111111111110",
										"1111111111111101",
										"1111111111111101",
										"1111111111111101",
										"1111111111111101",
										"1111111111111101",
										"1111111111111111",
										"1111111111111111",
										"0000000000000000",
										"0000000000000001",
										"0000000000000001",
										"0000000000000011",
										"0000000000000100",
										"0000000000000101",
										"0000000000000110",
										"0000000000000110",
										"0000000000000110",
										"0000000000000101",
										"0000000000000100",
										"0000000000000100",
										"0000000000000100",
										"0000000000000011",
										"0000000000000011",
										"0000000000000100",
										"0000000000000100",
										"0000000000000101",
										"0000000000000110",
										"0000000000000110",
										"0000000000000101",
										"0000000000000100",
										"0000000000000011",
										"0000000000000010",
										"0000000000000011",
										"0000000000000100",
										"0000000000000100",
										"0000000000000101",
										"0000000000000110",
										"0000000000000110",
										"0000000000000111",
										"0000000000000111",
										"0000000000000110",
										"0000000000000101",
										"0000000000000011",
										"0000000000000001",
										"0000000000000001",
										"0000000000000010",
										"0000000000000010",
										"0000000000000011",
										"0000000000000011",
										"0000000000000100",
										"0000000000000111",
										"0000000000001001",
										"0000000000001011",
										"0000000000001100",
										"0000000000001011",
										"0000000000001010",
										"0000000000001001",
										"0000000000001000",
										"0000000000000111",
										"0000000000000101",
										"0000000000000100",
										"0000000000000011",
										"0000000000000011",
										"0000000000000011",
										"0000000000000001",
										"0000000000000000",
										"0000000000000000",
										"0000000000000010",
										"0000000000000101",
										"0000000000000101",
										"0000000000000101",
										"0000000000000011",
										"0000000000000001",
										"0000000000000010",
										"0000000000000011",
										"0000000000000011",
										"0000000000000010",
										"0000000000000010",
										"0000000000000000",
										"0000000000000000",
										"0000000000000001",
										"0000000000000000",
										"0000000000000001",
										"0000000000000010",
										"0000000000000010",
										"0000000000000010",
										"0000000000000010",
										"0000000000000001",
										"0000000000000010",
										"0000000000000011",
										"0000000000000011",
										"0000000000000100",
										"0000000000000100",
										"0000000000000011",
										"0000000000000011",
										"0000000000000011",
										"0000000000000010",
										"0000000000000010",
										"0000000000000010",
										"0000000000000001",
										"0000000000000000",
										"0000000000000001",
										"0000000000000000",
										"0000000000000000",
										"0000000000000010",
										"0000000000000010",
										"0000000000000010",
										"0000000000000010",
										"0000000000000000",
										"1111111111111110",
										"1111111111111110",
										"1111111111111111",
										"0000000000000001",
										"0000000000000011",
										"0000000000000011",
										"0000000000000011",
										"0000000000000100",
										"0000000000000100",
										"0000000000000101",
										"0000000000000101",
										"0000000000000010",
										"0000000000000000",
										"0000000000000000",
										"0000000000000000",
										"0000000000000001",
										"0000000000000010",
										"0000000000000001",
										"0000000000000001",
										"0000000000000010",
										"0000000000000001",
										"0000000000000001",
										"0000000000000001",
										"0000000000000010",
										"0000000000000011",
										"0000000000000100",
										"0000000000000100",
										"0000000000000010",
										"0000000000000011",
										"0000000000000011",
										"0000000000000001",
										"0000000000000010",
										"0000000000000010",
										"0000000000000010",
										"0000000000000100",
										"0000000000000011",
										"0000000000000001",
										"0000000000000001",
										"0000000000000000",
										"0000000000000000",
										"0000000000000010",
										"0000000000000010",
										"0000000000000010",
										"0000000000000010",
										"0000000000000001",
										"0000000000000001",
										"0000000000000010",
										"0000000000000001",
										"0000000000000001",
										"0000000000000001",
										"0000000000000001",
										"0000000000000100",
										"0000000000000111",
										"0000000000000111",
										"0000000000000110",
										"0000000000000110",
										"0000000000000101",
										"0000000000000101",
										"0000000000000110",
										"0000000000000110",
										"0000000000000110",
										"0000000000000111",
										"0000000000000111",
										"0000000000000110",
										"0000000000000110",
										"0000000000000110",
										"0000000000000111",
										"0000000000000111",
										"0000000000000110",
										"0000000000000101",
										"0000000000000101",
										"0000000000000100",
										"0000000000000100",
										"0000000000000100",
										"0000000000000010",
										"0000000000000010",
										"0000000000000001",
										"0000000000000000",
										"0000000000000001",
										"0000000000000001",
										"0000000000000010",
										"0000000000000011",
										"0000000000000001",
										"0000000000000001",
										"0000000000000001",
										"0000000000000001",
										"0000000000000010",
										"0000000000000011",
										"0000000000000100",
										"0000000000000101",
										"0000000000000110",
										"0000000000000110",
										"0000000000000101",
										"0000000000000100",
										"0000000000000011",
										"0000000000000011",
										"0000000000000100",
										"0000000000000101",
										"0000000000000111",
										"0000000000001000",
										"0000000000001000",
										"0000000000000111",
										"0000000000000100",
										"0000000000000001",
										"1111111111111111",
										"1111111111111111",
										"0000000000000001",
										"0000000000000100",
										"0000000000000110",
										"0000000000000110",
										"0000000000000101",
										"0000000000000100",
										"0000000000000100",
										"0000000000000100",
										"0000000000000101",
										"0000000000000101",
										"0000000000000011",
										"0000000000000001",
										"0000000000000000",
										"0000000000000010",
										"0000000000000011",
										"0000000000000100",
										"0000000000000110",
										"0000000000000100",
										"0000000000000011",
										"0000000000000100",
										"0000000000000011",
										"0000000000000010",
										"0000000000000010",
										"0000000000000010",
										"0000000000000010",
										"0000000000000011",
										"0000000000000100",
										"0000000000000101",
										"0000000000000110",
										"0000000000000101",
										"0000000000000101",
										"0000000000000110",
										"0000000000000110",
										"0000000000000111",
										"0000000000001001",
										"0000000000000110",
										"0000000000000100",
										"0000000000000100",
										"0000000000000010",
										"0000000000000010",
										"0000000000000011",
										"0000000000000011",
										"0000000000000011",
										"0000000000000100",
										"0000000000000100",
										"0000000000000100",
										"0000000000000011",
										"0000000000000011",
										"0000000000000010",
										"0000000000000010",
										"0000000000000011",
										"0000000000000011",
										"0000000000000100",
										"0000000000000100",
										"0000000000000100",
										"0000000000000011",
										"0000000000000001",
										"0000000000000000",
										"0000000000000000",
										"0000000000000001",
										"0000000000000011",
										"0000000000000100",
										"0000000000000011",
										"0000000000000010",
										"0000000000000001",
										"0000000000000000",
										"0000000000000001",
										"0000000000000001",
										"0000000000000000",
										"0000000000000000",
										"1111111111111111",
										"1111111111111110",
										"1111111111111111",
										"0000000000000000",
										"0000000000000001",
										"0000000000000011",
										"0000000000000010",
										"0000000000000001",
										"0000000000000001",
										"0000000000000001",
										"0000000000000011",
										"0000000000000011",
										"0000000000000010",
										"0000000000000010",
										"0000000000000001",
										"0000000000000001",
										"0000000000000010",
										"0000000000000010",
										"0000000000000100",
										"0000000000000101",
										"0000000000000100",
										"0000000000000011",
										"0000000000000011",
										"0000000000000100",
										"0000000000000101",
										"0000000000000110",
										"0000000000000101",
										"0000000000000100",
										"0000000000000011",
										"0000000000000011",
										"0000000000000100",
										"0000000000000101",
										"0000000000000101",
										"0000000000000101",
										"0000000000000110",
										"0000000000000101",
										"0000000000000101",
										"0000000000000110",
										"0000000000000100",
										"0000000000000100",
										"0000000000000110",
										"0000000000000100",
										"0000000000000010",
										"0000000000000010",
										"0000000000000001",
										"0000000000000010",
										"0000000000000101",
										"0000000000000101",
										"0000000000000100",
										"0000000000000100",
										"0000000000000011",
										"0000000000000011",
										"0000000000000100",
										"0000000000000011",
										"0000000000000010",
										"0000000000000010",
										"0000000000000000",
										"1111111111111111",
										"0000000000000001",
										"0000000000000001",
										"0000000000000010",
										"0000000000000101",
										"0000000000000110",
										"0000000000000111",
										"0000000000000111",
										"0000000000000111",
										"0000000000000110",
										"0000000000000101",
										"0000000000000110",
										"0000000000000101",
										"0000000000000100",
										"0000000000000100",
										"0000000000000100",
										"0000000000000011",
										"0000000000000010",
										"0000000000000010",
										"0000000000000010",
										"0000000000000011",
										"0000000000000011",
										"0000000000000010",
										"0000000000000010",
										"0000000000000001",
										"0000000000000001",
										"0000000000000001",
										"0000000000000000",
										"0000000000000001",
										"0000000000000011",
										"0000000000000110",
										"0000000000000110",
										"0000000000000101",
										"0000000000000101",
										"0000000000000010",
										"0000000000000010",
										"0000000000000010",
										"0000000000000000",
										"0000000000000000",
										"0000000000000001",
										"0000000000000001",
										"0000000000000001",
										"0000000000000010",
										"0000000000000010",
										"0000000000000100",
										"0000000000000110",
										"0000000000000110",
										"0000000000000110",
										"0000000000000101",
										"0000000000000011",
										"0000000000000011",
										"0000000000000101",
										"0000000000000110",
										"0000000000000111",
										"0000000000000111",
										"0000000000000101",
										"0000000000000011",
										"0000000000000011",
										"0000000000000010",
										"0000000000000001",
										"0000000000000010",
										"0000000000000001",
										"0000000000000001",
										"0000000000000010",
										"0000000000000010",
										"0000000000000010",
										"0000000000000010",
										"0000000000000001",
										"0000000000000000",
										"0000000000000000",
										"0000000000000000",
										"0000000000000001",
										"0000000000000010",
										"0000000000000010",
										"0000000000000011",
										"0000000000000100",
										"0000000000000100",
										"0000000000000100",
										"0000000000000101",
										"0000000000000101",
										"0000000000000101",
										"0000000000000110",
										"0000000000000101",
										"0000000000000100",
										"0000000000000100",
										"0000000000000100",
										"0000000000000101",
										"0000000000000110",
										"0000000000000110",
										"0000000000000110",
										"0000000000000100",
										"0000000000000011",
										"0000000000000011",
										"0000000000000010",
										"0000000000000001",
										"0000000000000000",
										"0000000000000000",
										"0000000000000000",
										"0000000000000010",
										"0000000000000011",
										"0000000000000011",
										"0000000000000101",
										"0000000000000101",
										"0000000000000101",
										"0000000000000100",
										"0000000000000001",
										"0000000000000000",
										"1111111111111111",
										"1111111111111111",
										"0000000000000001",
										"0000000000000000",
										"0000000000000000",
										"0000000000000001",
										"0000000000000001",
										"0000000000000010",
										"0000000000000010",
										"0000000000000001",
										"0000000000000001",
										"0000000000000010",
										"0000000000000100",
										"0000000000000110",
										"0000000000000110",
										"0000000000000101",
										"0000000000000011",
										"0000000000000011",
										"0000000000000011",
										"0000000000000101",
										"0000000000000110",
										"0000000000000100",
										"0000000000000011",
										"0000000000000010",
										"0000000000000001",
										"0000000000000010",
										"0000000000000011",
										"0000000000000011",
										"0000000000000011",
										"0000000000000011",
										"0000000000000011",
										"0000000000000011",
										"0000000000000011",
										"0000000000000010",
										"0000000000000001",
										"0000000000000001",
										"0000000000000011",
										"0000000000000100",
										"0000000000000110",
										"0000000000000110",
										"0000000000000110",
										"0000000000000110",
										"0000000000000110",
										"0000000000000111",
										"0000000000000110",
										"0000000000000111",
										"0000000000001000",
										"0000000000000111",
										"0000000000000111",
										"0000000000000111",
										"0000000000000100",
										"0000000000000011",
										"0000000000000100",
										"0000000000000100",
										"0000000000000101",
										"0000000000000111",
										"0000000000000111",
										"0000000000000110",
										"0000000000000110",
										"0000000000000110",
										"0000000000000101",
										"0000000000000101",
										"0000000000000111",
										"0000000000000111",
										"0000000000000111",
										"0000000000000111",
										"0000000000000101",
										"0000000000000011",
										"0000000000000010",
										"0000000000000010",
										"0000000000000011",
										"0000000000000101",
										"0000000000000101",
										"0000000000000011",
										"0000000000000001",
										"0000000000000000",
										"0000000000000010",
										"0000000000000110",
										"0000000000000110",
										"0000000000000101",
										"0000000000000101",
										"0000000000000100",
										"0000000000000110",
										"0000000000000111",
										"0000000000000100",
										"0000000000000001",
										"0000000000000000",
										"0000000000000001",
										"0000000000000011",
										"0000000000000101",
										"0000000000000101",
										"0000000000000011",
										"0000000000000011",
										"0000000000000011",
										"0000000000000001",
										"0000000000000001",
										"0000000000000001",
										"0000000000000000",
										"0000000000000000",
										"0000000000000001",
										"0000000000000001",
										"0000000000000001",
										"0000000000000001",
										"1111111111111111",
										"1111111111111111",
										"0000000000000001",
										"0000000000000010",
										"0000000000000011",
										"0000000000000100",
										"0000000000000010",
										"0000000000000010",
										"0000000000000100",
										"0000000000000011",
										"0000000000000011",
										"0000000000000100",
										"0000000000000011",
										"0000000000000101",
										"0000000000000111",
										"0000000000000111",
										"0000000000000110",
										"0000000000000100",
										"0000000000000011",
										"0000000000000010",
										"0000000000000010",
										"0000000000000001",
										"0000000000000001",
										"0000000000000011",
										"0000000000000101",
										"0000000000000101",
										"0000000000000100",
										"0000000000000011",
										"0000000000000001",
										"0000000000000001",
										"0000000000000010",
										"0000000000000001",
										"0000000000000001",
										"0000000000000011",
										"0000000000000010",
										"0000000000000001",
										"0000000000000001",
										"0000000000000000",
										"0000000000000001",
										"0000000000000011",
										"0000000000000011",
										"0000000000000010",
										"0000000000000010",
										"0000000000000010",
										"0000000000000010",
										"0000000000000011",
										"0000000000000100",
										"0000000000000100",
										"0000000000000110",
										"0000000000000110",
										"0000000000000011",
										"0000000000000010",
										"0000000000000001",
										"0000000000000001",
										"0000000000000100",
										"0000000000000101",
										"0000000000000100",
										"0000000000000100",
										"0000000000000011",
										"0000000000000011",
										"0000000000000100",
										"0000000000000011",
										"0000000000000011",
										"0000000000000011",
										"0000000000000010",
										"0000000000000001",
										"0000000000000010"
										);
	
	
	begin
		
		-- inital reset of the filter
		rst_l <= '0';
		wait until clk'event and clk='1';
		rst_l <= '1'; 
		
		-- loop over all the samples
		for i in 0 to SAMPLES-1 loop	
			
			sample <= input(i);
			expected <= expected_out(i);
			
			
			wait until clk'event and clk='1'; 
			
			-- If the actual output and the expected output
			-- mismatch, raise an asserion
			assert (output = expected)
			report "Mismatch for index i = " & integer'image(i)
			severity error;
			
		end loop;	 
		
		enable <= '0';
		end process;

end TB_Arch;

