library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity ddfs_lut_4096 is
  port (
    address : in  std_logic_vector(11 downto 0);
    dds_out : out std_logic_vector(5 downto 0) 
  );
end ddfs_lut_4096;

architecture rtl of ddfs_lut_4096 is
type LUT_t is array (natural range 0 to 4095) of integer;
constant LUT: LUT_t := (
    0 => 0,
    1 => 0,
    2 => 0,
    3 => 0,
    4 => 0,
    5 => 0,
    6 => 0,
    7 => 0,
    8 => 0,
    9 => 0,
    10 => 0,
    11 => 0,
    12 => 0,
    13 => 0,
    14 => 0,
    15 => 0,
    16 => 0,
    17 => 0,
    18 => 0,
    19 => 0,
    20 => 0,
    21 => 0,
    22 => 1,
    23 => 1,
    24 => 1,
    25 => 1,
    26 => 1,
    27 => 1,
    28 => 1,
    29 => 1,
    30 => 1,
    31 => 1,
    32 => 1,
    33 => 1,
    34 => 1,
    35 => 1,
    36 => 1,
    37 => 1,
    38 => 1,
    39 => 1,
    40 => 1,
    41 => 1,
    42 => 1,
    43 => 2,
    44 => 2,
    45 => 2,
    46 => 2,
    47 => 2,
    48 => 2,
    49 => 2,
    50 => 2,
    51 => 2,
    52 => 2,
    53 => 2,
    54 => 2,
    55 => 2,
    56 => 2,
    57 => 2,
    58 => 2,
    59 => 2,
    60 => 2,
    61 => 2,
    62 => 2,
    63 => 2,
    64 => 3,
    65 => 3,
    66 => 3,
    67 => 3,
    68 => 3,
    69 => 3,
    70 => 3,
    71 => 3,
    72 => 3,
    73 => 3,
    74 => 3,
    75 => 3,
    76 => 3,
    77 => 3,
    78 => 3,
    79 => 3,
    80 => 3,
    81 => 3,
    82 => 3,
    83 => 3,
    84 => 3,
    85 => 4,
    86 => 4,
    87 => 4,
    88 => 4,
    89 => 4,
    90 => 4,
    91 => 4,
    92 => 4,
    93 => 4,
    94 => 4,
    95 => 4,
    96 => 4,
    97 => 4,
    98 => 4,
    99 => 4,
    100 => 4,
    101 => 4,
    102 => 4,
    103 => 4,
    104 => 4,
    105 => 4,
    106 => 5,
    107 => 5,
    108 => 5,
    109 => 5,
    110 => 5,
    111 => 5,
    112 => 5,
    113 => 5,
    114 => 5,
    115 => 5,
    116 => 5,
    117 => 5,
    118 => 5,
    119 => 5,
    120 => 5,
    121 => 5,
    122 => 5,
    123 => 5,
    124 => 5,
    125 => 5,
    126 => 5,
    127 => 6,
    128 => 6,
    129 => 6,
    130 => 6,
    131 => 6,
    132 => 6,
    133 => 6,
    134 => 6,
    135 => 6,
    136 => 6,
    137 => 6,
    138 => 6,
    139 => 6,
    140 => 6,
    141 => 6,
    142 => 6,
    143 => 6,
    144 => 6,
    145 => 6,
    146 => 6,
    147 => 6,
    148 => 6,
    149 => 7,
    150 => 7,
    151 => 7,
    152 => 7,
    153 => 7,
    154 => 7,
    155 => 7,
    156 => 7,
    157 => 7,
    158 => 7,
    159 => 7,
    160 => 7,
    161 => 7,
    162 => 7,
    163 => 7,
    164 => 7,
    165 => 7,
    166 => 7,
    167 => 7,
    168 => 7,
    169 => 7,
    170 => 7,
    171 => 8,
    172 => 8,
    173 => 8,
    174 => 8,
    175 => 8,
    176 => 8,
    177 => 8,
    178 => 8,
    179 => 8,
    180 => 8,
    181 => 8,
    182 => 8,
    183 => 8,
    184 => 8,
    185 => 8,
    186 => 8,
    187 => 8,
    188 => 8,
    189 => 8,
    190 => 8,
    191 => 8,
    192 => 8,
    193 => 9,
    194 => 9,
    195 => 9,
    196 => 9,
    197 => 9,
    198 => 9,
    199 => 9,
    200 => 9,
    201 => 9,
    202 => 9,
    203 => 9,
    204 => 9,
    205 => 9,
    206 => 9,
    207 => 9,
    208 => 9,
    209 => 9,
    210 => 9,
    211 => 9,
    212 => 9,
    213 => 9,
    214 => 9,
    215 => 10,
    216 => 10,
    217 => 10,
    218 => 10,
    219 => 10,
    220 => 10,
    221 => 10,
    222 => 10,
    223 => 10,
    224 => 10,
    225 => 10,
    226 => 10,
    227 => 10,
    228 => 10,
    229 => 10,
    230 => 10,
    231 => 10,
    232 => 10,
    233 => 10,
    234 => 10,
    235 => 10,
    236 => 10,
    237 => 11,
    238 => 11,
    239 => 11,
    240 => 11,
    241 => 11,
    242 => 11,
    243 => 11,
    244 => 11,
    245 => 11,
    246 => 11,
    247 => 11,
    248 => 11,
    249 => 11,
    250 => 11,
    251 => 11,
    252 => 11,
    253 => 11,
    254 => 11,
    255 => 11,
    256 => 11,
    257 => 11,
    258 => 11,
    259 => 11,
    260 => 12,
    261 => 12,
    262 => 12,
    263 => 12,
    264 => 12,
    265 => 12,
    266 => 12,
    267 => 12,
    268 => 12,
    269 => 12,
    270 => 12,
    271 => 12,
    272 => 12,
    273 => 12,
    274 => 12,
    275 => 12,
    276 => 12,
    277 => 12,
    278 => 12,
    279 => 12,
    280 => 12,
    281 => 12,
    282 => 12,
    283 => 13,
    284 => 13,
    285 => 13,
    286 => 13,
    287 => 13,
    288 => 13,
    289 => 13,
    290 => 13,
    291 => 13,
    292 => 13,
    293 => 13,
    294 => 13,
    295 => 13,
    296 => 13,
    297 => 13,
    298 => 13,
    299 => 13,
    300 => 13,
    301 => 13,
    302 => 13,
    303 => 13,
    304 => 13,
    305 => 13,
    306 => 14,
    307 => 14,
    308 => 14,
    309 => 14,
    310 => 14,
    311 => 14,
    312 => 14,
    313 => 14,
    314 => 14,
    315 => 14,
    316 => 14,
    317 => 14,
    318 => 14,
    319 => 14,
    320 => 14,
    321 => 14,
    322 => 14,
    323 => 14,
    324 => 14,
    325 => 14,
    326 => 14,
    327 => 14,
    328 => 14,
    329 => 14,
    330 => 15,
    331 => 15,
    332 => 15,
    333 => 15,
    334 => 15,
    335 => 15,
    336 => 15,
    337 => 15,
    338 => 15,
    339 => 15,
    340 => 15,
    341 => 15,
    342 => 15,
    343 => 15,
    344 => 15,
    345 => 15,
    346 => 15,
    347 => 15,
    348 => 15,
    349 => 15,
    350 => 15,
    351 => 15,
    352 => 15,
    353 => 15,
    354 => 16,
    355 => 16,
    356 => 16,
    357 => 16,
    358 => 16,
    359 => 16,
    360 => 16,
    361 => 16,
    362 => 16,
    363 => 16,
    364 => 16,
    365 => 16,
    366 => 16,
    367 => 16,
    368 => 16,
    369 => 16,
    370 => 16,
    371 => 16,
    372 => 16,
    373 => 16,
    374 => 16,
    375 => 16,
    376 => 16,
    377 => 16,
    378 => 16,
    379 => 17,
    380 => 17,
    381 => 17,
    382 => 17,
    383 => 17,
    384 => 17,
    385 => 17,
    386 => 17,
    387 => 17,
    388 => 17,
    389 => 17,
    390 => 17,
    391 => 17,
    392 => 17,
    393 => 17,
    394 => 17,
    395 => 17,
    396 => 17,
    397 => 17,
    398 => 17,
    399 => 17,
    400 => 17,
    401 => 17,
    402 => 17,
    403 => 17,
    404 => 18,
    405 => 18,
    406 => 18,
    407 => 18,
    408 => 18,
    409 => 18,
    410 => 18,
    411 => 18,
    412 => 18,
    413 => 18,
    414 => 18,
    415 => 18,
    416 => 18,
    417 => 18,
    418 => 18,
    419 => 18,
    420 => 18,
    421 => 18,
    422 => 18,
    423 => 18,
    424 => 18,
    425 => 18,
    426 => 18,
    427 => 18,
    428 => 18,
    429 => 18,
    430 => 18,
    431 => 19,
    432 => 19,
    433 => 19,
    434 => 19,
    435 => 19,
    436 => 19,
    437 => 19,
    438 => 19,
    439 => 19,
    440 => 19,
    441 => 19,
    442 => 19,
    443 => 19,
    444 => 19,
    445 => 19,
    446 => 19,
    447 => 19,
    448 => 19,
    449 => 19,
    450 => 19,
    451 => 19,
    452 => 19,
    453 => 19,
    454 => 19,
    455 => 19,
    456 => 19,
    457 => 19,
    458 => 20,
    459 => 20,
    460 => 20,
    461 => 20,
    462 => 20,
    463 => 20,
    464 => 20,
    465 => 20,
    466 => 20,
    467 => 20,
    468 => 20,
    469 => 20,
    470 => 20,
    471 => 20,
    472 => 20,
    473 => 20,
    474 => 20,
    475 => 20,
    476 => 20,
    477 => 20,
    478 => 20,
    479 => 20,
    480 => 20,
    481 => 20,
    482 => 20,
    483 => 20,
    484 => 20,
    485 => 20,
    486 => 21,
    487 => 21,
    488 => 21,
    489 => 21,
    490 => 21,
    491 => 21,
    492 => 21,
    493 => 21,
    494 => 21,
    495 => 21,
    496 => 21,
    497 => 21,
    498 => 21,
    499 => 21,
    500 => 21,
    501 => 21,
    502 => 21,
    503 => 21,
    504 => 21,
    505 => 21,
    506 => 21,
    507 => 21,
    508 => 21,
    509 => 21,
    510 => 21,
    511 => 21,
    512 => 21,
    513 => 21,
    514 => 21,
    515 => 22,
    516 => 22,
    517 => 22,
    518 => 22,
    519 => 22,
    520 => 22,
    521 => 22,
    522 => 22,
    523 => 22,
    524 => 22,
    525 => 22,
    526 => 22,
    527 => 22,
    528 => 22,
    529 => 22,
    530 => 22,
    531 => 22,
    532 => 22,
    533 => 22,
    534 => 22,
    535 => 22,
    536 => 22,
    537 => 22,
    538 => 22,
    539 => 22,
    540 => 22,
    541 => 22,
    542 => 22,
    543 => 22,
    544 => 22,
    545 => 23,
    546 => 23,
    547 => 23,
    548 => 23,
    549 => 23,
    550 => 23,
    551 => 23,
    552 => 23,
    553 => 23,
    554 => 23,
    555 => 23,
    556 => 23,
    557 => 23,
    558 => 23,
    559 => 23,
    560 => 23,
    561 => 23,
    562 => 23,
    563 => 23,
    564 => 23,
    565 => 23,
    566 => 23,
    567 => 23,
    568 => 23,
    569 => 23,
    570 => 23,
    571 => 23,
    572 => 23,
    573 => 23,
    574 => 23,
    575 => 23,
    576 => 23,
    577 => 23,
    578 => 24,
    579 => 24,
    580 => 24,
    581 => 24,
    582 => 24,
    583 => 24,
    584 => 24,
    585 => 24,
    586 => 24,
    587 => 24,
    588 => 24,
    589 => 24,
    590 => 24,
    591 => 24,
    592 => 24,
    593 => 24,
    594 => 24,
    595 => 24,
    596 => 24,
    597 => 24,
    598 => 24,
    599 => 24,
    600 => 24,
    601 => 24,
    602 => 24,
    603 => 24,
    604 => 24,
    605 => 24,
    606 => 24,
    607 => 24,
    608 => 24,
    609 => 24,
    610 => 24,
    611 => 24,
    612 => 25,
    613 => 25,
    614 => 25,
    615 => 25,
    616 => 25,
    617 => 25,
    618 => 25,
    619 => 25,
    620 => 25,
    621 => 25,
    622 => 25,
    623 => 25,
    624 => 25,
    625 => 25,
    626 => 25,
    627 => 25,
    628 => 25,
    629 => 25,
    630 => 25,
    631 => 25,
    632 => 25,
    633 => 25,
    634 => 25,
    635 => 25,
    636 => 25,
    637 => 25,
    638 => 25,
    639 => 25,
    640 => 25,
    641 => 25,
    642 => 25,
    643 => 25,
    644 => 25,
    645 => 25,
    646 => 25,
    647 => 25,
    648 => 25,
    649 => 26,
    650 => 26,
    651 => 26,
    652 => 26,
    653 => 26,
    654 => 26,
    655 => 26,
    656 => 26,
    657 => 26,
    658 => 26,
    659 => 26,
    660 => 26,
    661 => 26,
    662 => 26,
    663 => 26,
    664 => 26,
    665 => 26,
    666 => 26,
    667 => 26,
    668 => 26,
    669 => 26,
    670 => 26,
    671 => 26,
    672 => 26,
    673 => 26,
    674 => 26,
    675 => 26,
    676 => 26,
    677 => 26,
    678 => 26,
    679 => 26,
    680 => 26,
    681 => 26,
    682 => 26,
    683 => 26,
    684 => 26,
    685 => 26,
    686 => 26,
    687 => 26,
    688 => 26,
    689 => 26,
    690 => 27,
    691 => 27,
    692 => 27,
    693 => 27,
    694 => 27,
    695 => 27,
    696 => 27,
    697 => 27,
    698 => 27,
    699 => 27,
    700 => 27,
    701 => 27,
    702 => 27,
    703 => 27,
    704 => 27,
    705 => 27,
    706 => 27,
    707 => 27,
    708 => 27,
    709 => 27,
    710 => 27,
    711 => 27,
    712 => 27,
    713 => 27,
    714 => 27,
    715 => 27,
    716 => 27,
    717 => 27,
    718 => 27,
    719 => 27,
    720 => 27,
    721 => 27,
    722 => 27,
    723 => 27,
    724 => 27,
    725 => 27,
    726 => 27,
    727 => 27,
    728 => 27,
    729 => 27,
    730 => 27,
    731 => 27,
    732 => 27,
    733 => 27,
    734 => 27,
    735 => 28,
    736 => 28,
    737 => 28,
    738 => 28,
    739 => 28,
    740 => 28,
    741 => 28,
    742 => 28,
    743 => 28,
    744 => 28,
    745 => 28,
    746 => 28,
    747 => 28,
    748 => 28,
    749 => 28,
    750 => 28,
    751 => 28,
    752 => 28,
    753 => 28,
    754 => 28,
    755 => 28,
    756 => 28,
    757 => 28,
    758 => 28,
    759 => 28,
    760 => 28,
    761 => 28,
    762 => 28,
    763 => 28,
    764 => 28,
    765 => 28,
    766 => 28,
    767 => 28,
    768 => 28,
    769 => 28,
    770 => 28,
    771 => 28,
    772 => 28,
    773 => 28,
    774 => 28,
    775 => 28,
    776 => 28,
    777 => 28,
    778 => 28,
    779 => 28,
    780 => 28,
    781 => 28,
    782 => 28,
    783 => 28,
    784 => 28,
    785 => 28,
    786 => 28,
    787 => 28,
    788 => 28,
    789 => 29,
    790 => 29,
    791 => 29,
    792 => 29,
    793 => 29,
    794 => 29,
    795 => 29,
    796 => 29,
    797 => 29,
    798 => 29,
    799 => 29,
    800 => 29,
    801 => 29,
    802 => 29,
    803 => 29,
    804 => 29,
    805 => 29,
    806 => 29,
    807 => 29,
    808 => 29,
    809 => 29,
    810 => 29,
    811 => 29,
    812 => 29,
    813 => 29,
    814 => 29,
    815 => 29,
    816 => 29,
    817 => 29,
    818 => 29,
    819 => 29,
    820 => 29,
    821 => 29,
    822 => 29,
    823 => 29,
    824 => 29,
    825 => 29,
    826 => 29,
    827 => 29,
    828 => 29,
    829 => 29,
    830 => 29,
    831 => 29,
    832 => 29,
    833 => 29,
    834 => 29,
    835 => 29,
    836 => 29,
    837 => 29,
    838 => 29,
    839 => 29,
    840 => 29,
    841 => 29,
    842 => 29,
    843 => 29,
    844 => 29,
    845 => 29,
    846 => 29,
    847 => 29,
    848 => 29,
    849 => 29,
    850 => 29,
    851 => 29,
    852 => 29,
    853 => 29,
    854 => 29,
    855 => 29,
    856 => 29,
    857 => 29,
    858 => 30,
    859 => 30,
    860 => 30,
    861 => 30,
    862 => 30,
    863 => 30,
    864 => 30,
    865 => 30,
    866 => 30,
    867 => 30,
    868 => 30,
    869 => 30,
    870 => 30,
    871 => 30,
    872 => 30,
    873 => 30,
    874 => 30,
    875 => 30,
    876 => 30,
    877 => 30,
    878 => 30,
    879 => 30,
    880 => 30,
    881 => 30,
    882 => 30,
    883 => 30,
    884 => 30,
    885 => 30,
    886 => 30,
    887 => 30,
    888 => 30,
    889 => 30,
    890 => 30,
    891 => 30,
    892 => 30,
    893 => 30,
    894 => 30,
    895 => 30,
    896 => 30,
    897 => 30,
    898 => 30,
    899 => 30,
    900 => 30,
    901 => 30,
    902 => 30,
    903 => 30,
    904 => 30,
    905 => 30,
    906 => 30,
    907 => 30,
    908 => 30,
    909 => 30,
    910 => 30,
    911 => 30,
    912 => 30,
    913 => 30,
    914 => 30,
    915 => 30,
    916 => 30,
    917 => 30,
    918 => 30,
    919 => 30,
    920 => 30,
    921 => 30,
    922 => 30,
    923 => 30,
    924 => 30,
    925 => 30,
    926 => 30,
    927 => 30,
    928 => 30,
    929 => 30,
    930 => 30,
    931 => 30,
    932 => 30,
    933 => 30,
    934 => 30,
    935 => 30,
    936 => 30,
    937 => 30,
    938 => 30,
    939 => 30,
    940 => 30,
    941 => 30,
    942 => 30,
    943 => 30,
    944 => 30,
    945 => 30,
    946 => 30,
    947 => 30,
    948 => 30,
    949 => 30,
    950 => 30,
    951 => 30,
    952 => 30,
    953 => 30,
    954 => 30,
    955 => 30,
    956 => 30,
    957 => 30,
    958 => 30,
    959 => 30,
    960 => 30,
    961 => 30,
    962 => 30,
    963 => 30,
    964 => 30,
    965 => 30,
    966 => 30,
    967 => 30,
    968 => 30,
    969 => 30,
    970 => 30,
    971 => 30,
    972 => 30,
    973 => 30,
    974 => 30,
    975 => 30,
    976 => 30,
    977 => 30,
    978 => 30,
    979 => 30,
    980 => 30,
    981 => 30,
    982 => 30,
    983 => 30,
    984 => 30,
    985 => 30,
    986 => 30,
    987 => 30,
    988 => 30,
    989 => 30,
    990 => 30,
    991 => 30,
    992 => 30,
    993 => 30,
    994 => 30,
    995 => 30,
    996 => 30,
    997 => 30,
    998 => 30,
    999 => 30,
    1000 => 30,
    1001 => 30,
    1002 => 30,
    1003 => 30,
    1004 => 30,
    1005 => 30,
    1006 => 30,
    1007 => 30,
    1008 => 30,
    1009 => 30,
    1010 => 30,
    1011 => 30,
    1012 => 30,
    1013 => 30,
    1014 => 30,
    1015 => 30,
    1016 => 30,
    1017 => 30,
    1018 => 30,
    1019 => 30,
    1020 => 30,
    1021 => 30,
    1022 => 30,
    1023 => 30,
    1024 => 31,
    1025 => 30,
    1026 => 30,
    1027 => 30,
    1028 => 30,
    1029 => 30,
    1030 => 30,
    1031 => 30,
    1032 => 30,
    1033 => 30,
    1034 => 30,
    1035 => 30,
    1036 => 30,
    1037 => 30,
    1038 => 30,
    1039 => 30,
    1040 => 30,
    1041 => 30,
    1042 => 30,
    1043 => 30,
    1044 => 30,
    1045 => 30,
    1046 => 30,
    1047 => 30,
    1048 => 30,
    1049 => 30,
    1050 => 30,
    1051 => 30,
    1052 => 30,
    1053 => 30,
    1054 => 30,
    1055 => 30,
    1056 => 30,
    1057 => 30,
    1058 => 30,
    1059 => 30,
    1060 => 30,
    1061 => 30,
    1062 => 30,
    1063 => 30,
    1064 => 30,
    1065 => 30,
    1066 => 30,
    1067 => 30,
    1068 => 30,
    1069 => 30,
    1070 => 30,
    1071 => 30,
    1072 => 30,
    1073 => 30,
    1074 => 30,
    1075 => 30,
    1076 => 30,
    1077 => 30,
    1078 => 30,
    1079 => 30,
    1080 => 30,
    1081 => 30,
    1082 => 30,
    1083 => 30,
    1084 => 30,
    1085 => 30,
    1086 => 30,
    1087 => 30,
    1088 => 30,
    1089 => 30,
    1090 => 30,
    1091 => 30,
    1092 => 30,
    1093 => 30,
    1094 => 30,
    1095 => 30,
    1096 => 30,
    1097 => 30,
    1098 => 30,
    1099 => 30,
    1100 => 30,
    1101 => 30,
    1102 => 30,
    1103 => 30,
    1104 => 30,
    1105 => 30,
    1106 => 30,
    1107 => 30,
    1108 => 30,
    1109 => 30,
    1110 => 30,
    1111 => 30,
    1112 => 30,
    1113 => 30,
    1114 => 30,
    1115 => 30,
    1116 => 30,
    1117 => 30,
    1118 => 30,
    1119 => 30,
    1120 => 30,
    1121 => 30,
    1122 => 30,
    1123 => 30,
    1124 => 30,
    1125 => 30,
    1126 => 30,
    1127 => 30,
    1128 => 30,
    1129 => 30,
    1130 => 30,
    1131 => 30,
    1132 => 30,
    1133 => 30,
    1134 => 30,
    1135 => 30,
    1136 => 30,
    1137 => 30,
    1138 => 30,
    1139 => 30,
    1140 => 30,
    1141 => 30,
    1142 => 30,
    1143 => 30,
    1144 => 30,
    1145 => 30,
    1146 => 30,
    1147 => 30,
    1148 => 30,
    1149 => 30,
    1150 => 30,
    1151 => 30,
    1152 => 30,
    1153 => 30,
    1154 => 30,
    1155 => 30,
    1156 => 30,
    1157 => 30,
    1158 => 30,
    1159 => 30,
    1160 => 30,
    1161 => 30,
    1162 => 30,
    1163 => 30,
    1164 => 30,
    1165 => 30,
    1166 => 30,
    1167 => 30,
    1168 => 30,
    1169 => 30,
    1170 => 30,
    1171 => 30,
    1172 => 30,
    1173 => 30,
    1174 => 30,
    1175 => 30,
    1176 => 30,
    1177 => 30,
    1178 => 30,
    1179 => 30,
    1180 => 30,
    1181 => 30,
    1182 => 30,
    1183 => 30,
    1184 => 30,
    1185 => 30,
    1186 => 30,
    1187 => 30,
    1188 => 30,
    1189 => 30,
    1190 => 30,
    1191 => 29,
    1192 => 29,
    1193 => 29,
    1194 => 29,
    1195 => 29,
    1196 => 29,
    1197 => 29,
    1198 => 29,
    1199 => 29,
    1200 => 29,
    1201 => 29,
    1202 => 29,
    1203 => 29,
    1204 => 29,
    1205 => 29,
    1206 => 29,
    1207 => 29,
    1208 => 29,
    1209 => 29,
    1210 => 29,
    1211 => 29,
    1212 => 29,
    1213 => 29,
    1214 => 29,
    1215 => 29,
    1216 => 29,
    1217 => 29,
    1218 => 29,
    1219 => 29,
    1220 => 29,
    1221 => 29,
    1222 => 29,
    1223 => 29,
    1224 => 29,
    1225 => 29,
    1226 => 29,
    1227 => 29,
    1228 => 29,
    1229 => 29,
    1230 => 29,
    1231 => 29,
    1232 => 29,
    1233 => 29,
    1234 => 29,
    1235 => 29,
    1236 => 29,
    1237 => 29,
    1238 => 29,
    1239 => 29,
    1240 => 29,
    1241 => 29,
    1242 => 29,
    1243 => 29,
    1244 => 29,
    1245 => 29,
    1246 => 29,
    1247 => 29,
    1248 => 29,
    1249 => 29,
    1250 => 29,
    1251 => 29,
    1252 => 29,
    1253 => 29,
    1254 => 29,
    1255 => 29,
    1256 => 29,
    1257 => 29,
    1258 => 29,
    1259 => 29,
    1260 => 28,
    1261 => 28,
    1262 => 28,
    1263 => 28,
    1264 => 28,
    1265 => 28,
    1266 => 28,
    1267 => 28,
    1268 => 28,
    1269 => 28,
    1270 => 28,
    1271 => 28,
    1272 => 28,
    1273 => 28,
    1274 => 28,
    1275 => 28,
    1276 => 28,
    1277 => 28,
    1278 => 28,
    1279 => 28,
    1280 => 28,
    1281 => 28,
    1282 => 28,
    1283 => 28,
    1284 => 28,
    1285 => 28,
    1286 => 28,
    1287 => 28,
    1288 => 28,
    1289 => 28,
    1290 => 28,
    1291 => 28,
    1292 => 28,
    1293 => 28,
    1294 => 28,
    1295 => 28,
    1296 => 28,
    1297 => 28,
    1298 => 28,
    1299 => 28,
    1300 => 28,
    1301 => 28,
    1302 => 28,
    1303 => 28,
    1304 => 28,
    1305 => 28,
    1306 => 28,
    1307 => 28,
    1308 => 28,
    1309 => 28,
    1310 => 28,
    1311 => 28,
    1312 => 28,
    1313 => 28,
    1314 => 27,
    1315 => 27,
    1316 => 27,
    1317 => 27,
    1318 => 27,
    1319 => 27,
    1320 => 27,
    1321 => 27,
    1322 => 27,
    1323 => 27,
    1324 => 27,
    1325 => 27,
    1326 => 27,
    1327 => 27,
    1328 => 27,
    1329 => 27,
    1330 => 27,
    1331 => 27,
    1332 => 27,
    1333 => 27,
    1334 => 27,
    1335 => 27,
    1336 => 27,
    1337 => 27,
    1338 => 27,
    1339 => 27,
    1340 => 27,
    1341 => 27,
    1342 => 27,
    1343 => 27,
    1344 => 27,
    1345 => 27,
    1346 => 27,
    1347 => 27,
    1348 => 27,
    1349 => 27,
    1350 => 27,
    1351 => 27,
    1352 => 27,
    1353 => 27,
    1354 => 27,
    1355 => 27,
    1356 => 27,
    1357 => 27,
    1358 => 27,
    1359 => 26,
    1360 => 26,
    1361 => 26,
    1362 => 26,
    1363 => 26,
    1364 => 26,
    1365 => 26,
    1366 => 26,
    1367 => 26,
    1368 => 26,
    1369 => 26,
    1370 => 26,
    1371 => 26,
    1372 => 26,
    1373 => 26,
    1374 => 26,
    1375 => 26,
    1376 => 26,
    1377 => 26,
    1378 => 26,
    1379 => 26,
    1380 => 26,
    1381 => 26,
    1382 => 26,
    1383 => 26,
    1384 => 26,
    1385 => 26,
    1386 => 26,
    1387 => 26,
    1388 => 26,
    1389 => 26,
    1390 => 26,
    1391 => 26,
    1392 => 26,
    1393 => 26,
    1394 => 26,
    1395 => 26,
    1396 => 26,
    1397 => 26,
    1398 => 26,
    1399 => 26,
    1400 => 25,
    1401 => 25,
    1402 => 25,
    1403 => 25,
    1404 => 25,
    1405 => 25,
    1406 => 25,
    1407 => 25,
    1408 => 25,
    1409 => 25,
    1410 => 25,
    1411 => 25,
    1412 => 25,
    1413 => 25,
    1414 => 25,
    1415 => 25,
    1416 => 25,
    1417 => 25,
    1418 => 25,
    1419 => 25,
    1420 => 25,
    1421 => 25,
    1422 => 25,
    1423 => 25,
    1424 => 25,
    1425 => 25,
    1426 => 25,
    1427 => 25,
    1428 => 25,
    1429 => 25,
    1430 => 25,
    1431 => 25,
    1432 => 25,
    1433 => 25,
    1434 => 25,
    1435 => 25,
    1436 => 25,
    1437 => 24,
    1438 => 24,
    1439 => 24,
    1440 => 24,
    1441 => 24,
    1442 => 24,
    1443 => 24,
    1444 => 24,
    1445 => 24,
    1446 => 24,
    1447 => 24,
    1448 => 24,
    1449 => 24,
    1450 => 24,
    1451 => 24,
    1452 => 24,
    1453 => 24,
    1454 => 24,
    1455 => 24,
    1456 => 24,
    1457 => 24,
    1458 => 24,
    1459 => 24,
    1460 => 24,
    1461 => 24,
    1462 => 24,
    1463 => 24,
    1464 => 24,
    1465 => 24,
    1466 => 24,
    1467 => 24,
    1468 => 24,
    1469 => 24,
    1470 => 24,
    1471 => 23,
    1472 => 23,
    1473 => 23,
    1474 => 23,
    1475 => 23,
    1476 => 23,
    1477 => 23,
    1478 => 23,
    1479 => 23,
    1480 => 23,
    1481 => 23,
    1482 => 23,
    1483 => 23,
    1484 => 23,
    1485 => 23,
    1486 => 23,
    1487 => 23,
    1488 => 23,
    1489 => 23,
    1490 => 23,
    1491 => 23,
    1492 => 23,
    1493 => 23,
    1494 => 23,
    1495 => 23,
    1496 => 23,
    1497 => 23,
    1498 => 23,
    1499 => 23,
    1500 => 23,
    1501 => 23,
    1502 => 23,
    1503 => 23,
    1504 => 22,
    1505 => 22,
    1506 => 22,
    1507 => 22,
    1508 => 22,
    1509 => 22,
    1510 => 22,
    1511 => 22,
    1512 => 22,
    1513 => 22,
    1514 => 22,
    1515 => 22,
    1516 => 22,
    1517 => 22,
    1518 => 22,
    1519 => 22,
    1520 => 22,
    1521 => 22,
    1522 => 22,
    1523 => 22,
    1524 => 22,
    1525 => 22,
    1526 => 22,
    1527 => 22,
    1528 => 22,
    1529 => 22,
    1530 => 22,
    1531 => 22,
    1532 => 22,
    1533 => 22,
    1534 => 21,
    1535 => 21,
    1536 => 21,
    1537 => 21,
    1538 => 21,
    1539 => 21,
    1540 => 21,
    1541 => 21,
    1542 => 21,
    1543 => 21,
    1544 => 21,
    1545 => 21,
    1546 => 21,
    1547 => 21,
    1548 => 21,
    1549 => 21,
    1550 => 21,
    1551 => 21,
    1552 => 21,
    1553 => 21,
    1554 => 21,
    1555 => 21,
    1556 => 21,
    1557 => 21,
    1558 => 21,
    1559 => 21,
    1560 => 21,
    1561 => 21,
    1562 => 21,
    1563 => 20,
    1564 => 20,
    1565 => 20,
    1566 => 20,
    1567 => 20,
    1568 => 20,
    1569 => 20,
    1570 => 20,
    1571 => 20,
    1572 => 20,
    1573 => 20,
    1574 => 20,
    1575 => 20,
    1576 => 20,
    1577 => 20,
    1578 => 20,
    1579 => 20,
    1580 => 20,
    1581 => 20,
    1582 => 20,
    1583 => 20,
    1584 => 20,
    1585 => 20,
    1586 => 20,
    1587 => 20,
    1588 => 20,
    1589 => 20,
    1590 => 20,
    1591 => 19,
    1592 => 19,
    1593 => 19,
    1594 => 19,
    1595 => 19,
    1596 => 19,
    1597 => 19,
    1598 => 19,
    1599 => 19,
    1600 => 19,
    1601 => 19,
    1602 => 19,
    1603 => 19,
    1604 => 19,
    1605 => 19,
    1606 => 19,
    1607 => 19,
    1608 => 19,
    1609 => 19,
    1610 => 19,
    1611 => 19,
    1612 => 19,
    1613 => 19,
    1614 => 19,
    1615 => 19,
    1616 => 19,
    1617 => 19,
    1618 => 18,
    1619 => 18,
    1620 => 18,
    1621 => 18,
    1622 => 18,
    1623 => 18,
    1624 => 18,
    1625 => 18,
    1626 => 18,
    1627 => 18,
    1628 => 18,
    1629 => 18,
    1630 => 18,
    1631 => 18,
    1632 => 18,
    1633 => 18,
    1634 => 18,
    1635 => 18,
    1636 => 18,
    1637 => 18,
    1638 => 18,
    1639 => 18,
    1640 => 18,
    1641 => 18,
    1642 => 18,
    1643 => 18,
    1644 => 18,
    1645 => 17,
    1646 => 17,
    1647 => 17,
    1648 => 17,
    1649 => 17,
    1650 => 17,
    1651 => 17,
    1652 => 17,
    1653 => 17,
    1654 => 17,
    1655 => 17,
    1656 => 17,
    1657 => 17,
    1658 => 17,
    1659 => 17,
    1660 => 17,
    1661 => 17,
    1662 => 17,
    1663 => 17,
    1664 => 17,
    1665 => 17,
    1666 => 17,
    1667 => 17,
    1668 => 17,
    1669 => 17,
    1670 => 16,
    1671 => 16,
    1672 => 16,
    1673 => 16,
    1674 => 16,
    1675 => 16,
    1676 => 16,
    1677 => 16,
    1678 => 16,
    1679 => 16,
    1680 => 16,
    1681 => 16,
    1682 => 16,
    1683 => 16,
    1684 => 16,
    1685 => 16,
    1686 => 16,
    1687 => 16,
    1688 => 16,
    1689 => 16,
    1690 => 16,
    1691 => 16,
    1692 => 16,
    1693 => 16,
    1694 => 16,
    1695 => 15,
    1696 => 15,
    1697 => 15,
    1698 => 15,
    1699 => 15,
    1700 => 15,
    1701 => 15,
    1702 => 15,
    1703 => 15,
    1704 => 15,
    1705 => 15,
    1706 => 15,
    1707 => 15,
    1708 => 15,
    1709 => 15,
    1710 => 15,
    1711 => 15,
    1712 => 15,
    1713 => 15,
    1714 => 15,
    1715 => 15,
    1716 => 15,
    1717 => 15,
    1718 => 15,
    1719 => 14,
    1720 => 14,
    1721 => 14,
    1722 => 14,
    1723 => 14,
    1724 => 14,
    1725 => 14,
    1726 => 14,
    1727 => 14,
    1728 => 14,
    1729 => 14,
    1730 => 14,
    1731 => 14,
    1732 => 14,
    1733 => 14,
    1734 => 14,
    1735 => 14,
    1736 => 14,
    1737 => 14,
    1738 => 14,
    1739 => 14,
    1740 => 14,
    1741 => 14,
    1742 => 14,
    1743 => 13,
    1744 => 13,
    1745 => 13,
    1746 => 13,
    1747 => 13,
    1748 => 13,
    1749 => 13,
    1750 => 13,
    1751 => 13,
    1752 => 13,
    1753 => 13,
    1754 => 13,
    1755 => 13,
    1756 => 13,
    1757 => 13,
    1758 => 13,
    1759 => 13,
    1760 => 13,
    1761 => 13,
    1762 => 13,
    1763 => 13,
    1764 => 13,
    1765 => 13,
    1766 => 12,
    1767 => 12,
    1768 => 12,
    1769 => 12,
    1770 => 12,
    1771 => 12,
    1772 => 12,
    1773 => 12,
    1774 => 12,
    1775 => 12,
    1776 => 12,
    1777 => 12,
    1778 => 12,
    1779 => 12,
    1780 => 12,
    1781 => 12,
    1782 => 12,
    1783 => 12,
    1784 => 12,
    1785 => 12,
    1786 => 12,
    1787 => 12,
    1788 => 12,
    1789 => 11,
    1790 => 11,
    1791 => 11,
    1792 => 11,
    1793 => 11,
    1794 => 11,
    1795 => 11,
    1796 => 11,
    1797 => 11,
    1798 => 11,
    1799 => 11,
    1800 => 11,
    1801 => 11,
    1802 => 11,
    1803 => 11,
    1804 => 11,
    1805 => 11,
    1806 => 11,
    1807 => 11,
    1808 => 11,
    1809 => 11,
    1810 => 11,
    1811 => 11,
    1812 => 10,
    1813 => 10,
    1814 => 10,
    1815 => 10,
    1816 => 10,
    1817 => 10,
    1818 => 10,
    1819 => 10,
    1820 => 10,
    1821 => 10,
    1822 => 10,
    1823 => 10,
    1824 => 10,
    1825 => 10,
    1826 => 10,
    1827 => 10,
    1828 => 10,
    1829 => 10,
    1830 => 10,
    1831 => 10,
    1832 => 10,
    1833 => 10,
    1834 => 9,
    1835 => 9,
    1836 => 9,
    1837 => 9,
    1838 => 9,
    1839 => 9,
    1840 => 9,
    1841 => 9,
    1842 => 9,
    1843 => 9,
    1844 => 9,
    1845 => 9,
    1846 => 9,
    1847 => 9,
    1848 => 9,
    1849 => 9,
    1850 => 9,
    1851 => 9,
    1852 => 9,
    1853 => 9,
    1854 => 9,
    1855 => 9,
    1856 => 8,
    1857 => 8,
    1858 => 8,
    1859 => 8,
    1860 => 8,
    1861 => 8,
    1862 => 8,
    1863 => 8,
    1864 => 8,
    1865 => 8,
    1866 => 8,
    1867 => 8,
    1868 => 8,
    1869 => 8,
    1870 => 8,
    1871 => 8,
    1872 => 8,
    1873 => 8,
    1874 => 8,
    1875 => 8,
    1876 => 8,
    1877 => 8,
    1878 => 7,
    1879 => 7,
    1880 => 7,
    1881 => 7,
    1882 => 7,
    1883 => 7,
    1884 => 7,
    1885 => 7,
    1886 => 7,
    1887 => 7,
    1888 => 7,
    1889 => 7,
    1890 => 7,
    1891 => 7,
    1892 => 7,
    1893 => 7,
    1894 => 7,
    1895 => 7,
    1896 => 7,
    1897 => 7,
    1898 => 7,
    1899 => 7,
    1900 => 6,
    1901 => 6,
    1902 => 6,
    1903 => 6,
    1904 => 6,
    1905 => 6,
    1906 => 6,
    1907 => 6,
    1908 => 6,
    1909 => 6,
    1910 => 6,
    1911 => 6,
    1912 => 6,
    1913 => 6,
    1914 => 6,
    1915 => 6,
    1916 => 6,
    1917 => 6,
    1918 => 6,
    1919 => 6,
    1920 => 6,
    1921 => 6,
    1922 => 5,
    1923 => 5,
    1924 => 5,
    1925 => 5,
    1926 => 5,
    1927 => 5,
    1928 => 5,
    1929 => 5,
    1930 => 5,
    1931 => 5,
    1932 => 5,
    1933 => 5,
    1934 => 5,
    1935 => 5,
    1936 => 5,
    1937 => 5,
    1938 => 5,
    1939 => 5,
    1940 => 5,
    1941 => 5,
    1942 => 5,
    1943 => 4,
    1944 => 4,
    1945 => 4,
    1946 => 4,
    1947 => 4,
    1948 => 4,
    1949 => 4,
    1950 => 4,
    1951 => 4,
    1952 => 4,
    1953 => 4,
    1954 => 4,
    1955 => 4,
    1956 => 4,
    1957 => 4,
    1958 => 4,
    1959 => 4,
    1960 => 4,
    1961 => 4,
    1962 => 4,
    1963 => 4,
    1964 => 3,
    1965 => 3,
    1966 => 3,
    1967 => 3,
    1968 => 3,
    1969 => 3,
    1970 => 3,
    1971 => 3,
    1972 => 3,
    1973 => 3,
    1974 => 3,
    1975 => 3,
    1976 => 3,
    1977 => 3,
    1978 => 3,
    1979 => 3,
    1980 => 3,
    1981 => 3,
    1982 => 3,
    1983 => 3,
    1984 => 3,
    1985 => 2,
    1986 => 2,
    1987 => 2,
    1988 => 2,
    1989 => 2,
    1990 => 2,
    1991 => 2,
    1992 => 2,
    1993 => 2,
    1994 => 2,
    1995 => 2,
    1996 => 2,
    1997 => 2,
    1998 => 2,
    1999 => 2,
    2000 => 2,
    2001 => 2,
    2002 => 2,
    2003 => 2,
    2004 => 2,
    2005 => 2,
    2006 => 1,
    2007 => 1,
    2008 => 1,
    2009 => 1,
    2010 => 1,
    2011 => 1,
    2012 => 1,
    2013 => 1,
    2014 => 1,
    2015 => 1,
    2016 => 1,
    2017 => 1,
    2018 => 1,
    2019 => 1,
    2020 => 1,
    2021 => 1,
    2022 => 1,
    2023 => 1,
    2024 => 1,
    2025 => 1,
    2026 => 1,
    2027 => 0,
    2028 => 0,
    2029 => 0,
    2030 => 0,
    2031 => 0,
    2032 => 0,
    2033 => 0,
    2034 => 0,
    2035 => 0,
    2036 => 0,
    2037 => 0,
    2038 => 0,
    2039 => 0,
    2040 => 0,
    2041 => 0,
    2042 => 0,
    2043 => 0,
    2044 => 0,
    2045 => 0,
    2046 => 0,
    2047 => 0,
    2048 => 0,
    2049 => -1,
    2050 => -1,
    2051 => -1,
    2052 => -1,
    2053 => -1,
    2054 => -1,
    2055 => -1,
    2056 => -1,
    2057 => -1,
    2058 => -1,
    2059 => -1,
    2060 => -1,
    2061 => -1,
    2062 => -1,
    2063 => -1,
    2064 => -1,
    2065 => -1,
    2066 => -1,
    2067 => -1,
    2068 => -1,
    2069 => -1,
    2070 => -2,
    2071 => -2,
    2072 => -2,
    2073 => -2,
    2074 => -2,
    2075 => -2,
    2076 => -2,
    2077 => -2,
    2078 => -2,
    2079 => -2,
    2080 => -2,
    2081 => -2,
    2082 => -2,
    2083 => -2,
    2084 => -2,
    2085 => -2,
    2086 => -2,
    2087 => -2,
    2088 => -2,
    2089 => -2,
    2090 => -2,
    2091 => -3,
    2092 => -3,
    2093 => -3,
    2094 => -3,
    2095 => -3,
    2096 => -3,
    2097 => -3,
    2098 => -3,
    2099 => -3,
    2100 => -3,
    2101 => -3,
    2102 => -3,
    2103 => -3,
    2104 => -3,
    2105 => -3,
    2106 => -3,
    2107 => -3,
    2108 => -3,
    2109 => -3,
    2110 => -3,
    2111 => -3,
    2112 => -4,
    2113 => -4,
    2114 => -4,
    2115 => -4,
    2116 => -4,
    2117 => -4,
    2118 => -4,
    2119 => -4,
    2120 => -4,
    2121 => -4,
    2122 => -4,
    2123 => -4,
    2124 => -4,
    2125 => -4,
    2126 => -4,
    2127 => -4,
    2128 => -4,
    2129 => -4,
    2130 => -4,
    2131 => -4,
    2132 => -4,
    2133 => -5,
    2134 => -5,
    2135 => -5,
    2136 => -5,
    2137 => -5,
    2138 => -5,
    2139 => -5,
    2140 => -5,
    2141 => -5,
    2142 => -5,
    2143 => -5,
    2144 => -5,
    2145 => -5,
    2146 => -5,
    2147 => -5,
    2148 => -5,
    2149 => -5,
    2150 => -5,
    2151 => -5,
    2152 => -5,
    2153 => -5,
    2154 => -6,
    2155 => -6,
    2156 => -6,
    2157 => -6,
    2158 => -6,
    2159 => -6,
    2160 => -6,
    2161 => -6,
    2162 => -6,
    2163 => -6,
    2164 => -6,
    2165 => -6,
    2166 => -6,
    2167 => -6,
    2168 => -6,
    2169 => -6,
    2170 => -6,
    2171 => -6,
    2172 => -6,
    2173 => -6,
    2174 => -6,
    2175 => -7,
    2176 => -7,
    2177 => -7,
    2178 => -7,
    2179 => -7,
    2180 => -7,
    2181 => -7,
    2182 => -7,
    2183 => -7,
    2184 => -7,
    2185 => -7,
    2186 => -7,
    2187 => -7,
    2188 => -7,
    2189 => -7,
    2190 => -7,
    2191 => -7,
    2192 => -7,
    2193 => -7,
    2194 => -7,
    2195 => -7,
    2196 => -7,
    2197 => -8,
    2198 => -8,
    2199 => -8,
    2200 => -8,
    2201 => -8,
    2202 => -8,
    2203 => -8,
    2204 => -8,
    2205 => -8,
    2206 => -8,
    2207 => -8,
    2208 => -8,
    2209 => -8,
    2210 => -8,
    2211 => -8,
    2212 => -8,
    2213 => -8,
    2214 => -8,
    2215 => -8,
    2216 => -8,
    2217 => -8,
    2218 => -8,
    2219 => -9,
    2220 => -9,
    2221 => -9,
    2222 => -9,
    2223 => -9,
    2224 => -9,
    2225 => -9,
    2226 => -9,
    2227 => -9,
    2228 => -9,
    2229 => -9,
    2230 => -9,
    2231 => -9,
    2232 => -9,
    2233 => -9,
    2234 => -9,
    2235 => -9,
    2236 => -9,
    2237 => -9,
    2238 => -9,
    2239 => -9,
    2240 => -9,
    2241 => -10,
    2242 => -10,
    2243 => -10,
    2244 => -10,
    2245 => -10,
    2246 => -10,
    2247 => -10,
    2248 => -10,
    2249 => -10,
    2250 => -10,
    2251 => -10,
    2252 => -10,
    2253 => -10,
    2254 => -10,
    2255 => -10,
    2256 => -10,
    2257 => -10,
    2258 => -10,
    2259 => -10,
    2260 => -10,
    2261 => -10,
    2262 => -10,
    2263 => -11,
    2264 => -11,
    2265 => -11,
    2266 => -11,
    2267 => -11,
    2268 => -11,
    2269 => -11,
    2270 => -11,
    2271 => -11,
    2272 => -11,
    2273 => -11,
    2274 => -11,
    2275 => -11,
    2276 => -11,
    2277 => -11,
    2278 => -11,
    2279 => -11,
    2280 => -11,
    2281 => -11,
    2282 => -11,
    2283 => -11,
    2284 => -11,
    2285 => -12,
    2286 => -12,
    2287 => -12,
    2288 => -12,
    2289 => -12,
    2290 => -12,
    2291 => -12,
    2292 => -12,
    2293 => -12,
    2294 => -12,
    2295 => -12,
    2296 => -12,
    2297 => -12,
    2298 => -12,
    2299 => -12,
    2300 => -12,
    2301 => -12,
    2302 => -12,
    2303 => -12,
    2304 => -12,
    2305 => -12,
    2306 => -12,
    2307 => -12,
    2308 => -13,
    2309 => -13,
    2310 => -13,
    2311 => -13,
    2312 => -13,
    2313 => -13,
    2314 => -13,
    2315 => -13,
    2316 => -13,
    2317 => -13,
    2318 => -13,
    2319 => -13,
    2320 => -13,
    2321 => -13,
    2322 => -13,
    2323 => -13,
    2324 => -13,
    2325 => -13,
    2326 => -13,
    2327 => -13,
    2328 => -13,
    2329 => -13,
    2330 => -13,
    2331 => -14,
    2332 => -14,
    2333 => -14,
    2334 => -14,
    2335 => -14,
    2336 => -14,
    2337 => -14,
    2338 => -14,
    2339 => -14,
    2340 => -14,
    2341 => -14,
    2342 => -14,
    2343 => -14,
    2344 => -14,
    2345 => -14,
    2346 => -14,
    2347 => -14,
    2348 => -14,
    2349 => -14,
    2350 => -14,
    2351 => -14,
    2352 => -14,
    2353 => -14,
    2354 => -15,
    2355 => -15,
    2356 => -15,
    2357 => -15,
    2358 => -15,
    2359 => -15,
    2360 => -15,
    2361 => -15,
    2362 => -15,
    2363 => -15,
    2364 => -15,
    2365 => -15,
    2366 => -15,
    2367 => -15,
    2368 => -15,
    2369 => -15,
    2370 => -15,
    2371 => -15,
    2372 => -15,
    2373 => -15,
    2374 => -15,
    2375 => -15,
    2376 => -15,
    2377 => -15,
    2378 => -16,
    2379 => -16,
    2380 => -16,
    2381 => -16,
    2382 => -16,
    2383 => -16,
    2384 => -16,
    2385 => -16,
    2386 => -16,
    2387 => -16,
    2388 => -16,
    2389 => -16,
    2390 => -16,
    2391 => -16,
    2392 => -16,
    2393 => -16,
    2394 => -16,
    2395 => -16,
    2396 => -16,
    2397 => -16,
    2398 => -16,
    2399 => -16,
    2400 => -16,
    2401 => -16,
    2402 => -17,
    2403 => -17,
    2404 => -17,
    2405 => -17,
    2406 => -17,
    2407 => -17,
    2408 => -17,
    2409 => -17,
    2410 => -17,
    2411 => -17,
    2412 => -17,
    2413 => -17,
    2414 => -17,
    2415 => -17,
    2416 => -17,
    2417 => -17,
    2418 => -17,
    2419 => -17,
    2420 => -17,
    2421 => -17,
    2422 => -17,
    2423 => -17,
    2424 => -17,
    2425 => -17,
    2426 => -17,
    2427 => -18,
    2428 => -18,
    2429 => -18,
    2430 => -18,
    2431 => -18,
    2432 => -18,
    2433 => -18,
    2434 => -18,
    2435 => -18,
    2436 => -18,
    2437 => -18,
    2438 => -18,
    2439 => -18,
    2440 => -18,
    2441 => -18,
    2442 => -18,
    2443 => -18,
    2444 => -18,
    2445 => -18,
    2446 => -18,
    2447 => -18,
    2448 => -18,
    2449 => -18,
    2450 => -18,
    2451 => -18,
    2452 => -19,
    2453 => -19,
    2454 => -19,
    2455 => -19,
    2456 => -19,
    2457 => -19,
    2458 => -19,
    2459 => -19,
    2460 => -19,
    2461 => -19,
    2462 => -19,
    2463 => -19,
    2464 => -19,
    2465 => -19,
    2466 => -19,
    2467 => -19,
    2468 => -19,
    2469 => -19,
    2470 => -19,
    2471 => -19,
    2472 => -19,
    2473 => -19,
    2474 => -19,
    2475 => -19,
    2476 => -19,
    2477 => -19,
    2478 => -19,
    2479 => -20,
    2480 => -20,
    2481 => -20,
    2482 => -20,
    2483 => -20,
    2484 => -20,
    2485 => -20,
    2486 => -20,
    2487 => -20,
    2488 => -20,
    2489 => -20,
    2490 => -20,
    2491 => -20,
    2492 => -20,
    2493 => -20,
    2494 => -20,
    2495 => -20,
    2496 => -20,
    2497 => -20,
    2498 => -20,
    2499 => -20,
    2500 => -20,
    2501 => -20,
    2502 => -20,
    2503 => -20,
    2504 => -20,
    2505 => -20,
    2506 => -21,
    2507 => -21,
    2508 => -21,
    2509 => -21,
    2510 => -21,
    2511 => -21,
    2512 => -21,
    2513 => -21,
    2514 => -21,
    2515 => -21,
    2516 => -21,
    2517 => -21,
    2518 => -21,
    2519 => -21,
    2520 => -21,
    2521 => -21,
    2522 => -21,
    2523 => -21,
    2524 => -21,
    2525 => -21,
    2526 => -21,
    2527 => -21,
    2528 => -21,
    2529 => -21,
    2530 => -21,
    2531 => -21,
    2532 => -21,
    2533 => -21,
    2534 => -22,
    2535 => -22,
    2536 => -22,
    2537 => -22,
    2538 => -22,
    2539 => -22,
    2540 => -22,
    2541 => -22,
    2542 => -22,
    2543 => -22,
    2544 => -22,
    2545 => -22,
    2546 => -22,
    2547 => -22,
    2548 => -22,
    2549 => -22,
    2550 => -22,
    2551 => -22,
    2552 => -22,
    2553 => -22,
    2554 => -22,
    2555 => -22,
    2556 => -22,
    2557 => -22,
    2558 => -22,
    2559 => -22,
    2560 => -22,
    2561 => -22,
    2562 => -22,
    2563 => -23,
    2564 => -23,
    2565 => -23,
    2566 => -23,
    2567 => -23,
    2568 => -23,
    2569 => -23,
    2570 => -23,
    2571 => -23,
    2572 => -23,
    2573 => -23,
    2574 => -23,
    2575 => -23,
    2576 => -23,
    2577 => -23,
    2578 => -23,
    2579 => -23,
    2580 => -23,
    2581 => -23,
    2582 => -23,
    2583 => -23,
    2584 => -23,
    2585 => -23,
    2586 => -23,
    2587 => -23,
    2588 => -23,
    2589 => -23,
    2590 => -23,
    2591 => -23,
    2592 => -23,
    2593 => -24,
    2594 => -24,
    2595 => -24,
    2596 => -24,
    2597 => -24,
    2598 => -24,
    2599 => -24,
    2600 => -24,
    2601 => -24,
    2602 => -24,
    2603 => -24,
    2604 => -24,
    2605 => -24,
    2606 => -24,
    2607 => -24,
    2608 => -24,
    2609 => -24,
    2610 => -24,
    2611 => -24,
    2612 => -24,
    2613 => -24,
    2614 => -24,
    2615 => -24,
    2616 => -24,
    2617 => -24,
    2618 => -24,
    2619 => -24,
    2620 => -24,
    2621 => -24,
    2622 => -24,
    2623 => -24,
    2624 => -24,
    2625 => -24,
    2626 => -25,
    2627 => -25,
    2628 => -25,
    2629 => -25,
    2630 => -25,
    2631 => -25,
    2632 => -25,
    2633 => -25,
    2634 => -25,
    2635 => -25,
    2636 => -25,
    2637 => -25,
    2638 => -25,
    2639 => -25,
    2640 => -25,
    2641 => -25,
    2642 => -25,
    2643 => -25,
    2644 => -25,
    2645 => -25,
    2646 => -25,
    2647 => -25,
    2648 => -25,
    2649 => -25,
    2650 => -25,
    2651 => -25,
    2652 => -25,
    2653 => -25,
    2654 => -25,
    2655 => -25,
    2656 => -25,
    2657 => -25,
    2658 => -25,
    2659 => -25,
    2660 => -26,
    2661 => -26,
    2662 => -26,
    2663 => -26,
    2664 => -26,
    2665 => -26,
    2666 => -26,
    2667 => -26,
    2668 => -26,
    2669 => -26,
    2670 => -26,
    2671 => -26,
    2672 => -26,
    2673 => -26,
    2674 => -26,
    2675 => -26,
    2676 => -26,
    2677 => -26,
    2678 => -26,
    2679 => -26,
    2680 => -26,
    2681 => -26,
    2682 => -26,
    2683 => -26,
    2684 => -26,
    2685 => -26,
    2686 => -26,
    2687 => -26,
    2688 => -26,
    2689 => -26,
    2690 => -26,
    2691 => -26,
    2692 => -26,
    2693 => -26,
    2694 => -26,
    2695 => -26,
    2696 => -26,
    2697 => -27,
    2698 => -27,
    2699 => -27,
    2700 => -27,
    2701 => -27,
    2702 => -27,
    2703 => -27,
    2704 => -27,
    2705 => -27,
    2706 => -27,
    2707 => -27,
    2708 => -27,
    2709 => -27,
    2710 => -27,
    2711 => -27,
    2712 => -27,
    2713 => -27,
    2714 => -27,
    2715 => -27,
    2716 => -27,
    2717 => -27,
    2718 => -27,
    2719 => -27,
    2720 => -27,
    2721 => -27,
    2722 => -27,
    2723 => -27,
    2724 => -27,
    2725 => -27,
    2726 => -27,
    2727 => -27,
    2728 => -27,
    2729 => -27,
    2730 => -27,
    2731 => -27,
    2732 => -27,
    2733 => -27,
    2734 => -27,
    2735 => -27,
    2736 => -27,
    2737 => -27,
    2738 => -28,
    2739 => -28,
    2740 => -28,
    2741 => -28,
    2742 => -28,
    2743 => -28,
    2744 => -28,
    2745 => -28,
    2746 => -28,
    2747 => -28,
    2748 => -28,
    2749 => -28,
    2750 => -28,
    2751 => -28,
    2752 => -28,
    2753 => -28,
    2754 => -28,
    2755 => -28,
    2756 => -28,
    2757 => -28,
    2758 => -28,
    2759 => -28,
    2760 => -28,
    2761 => -28,
    2762 => -28,
    2763 => -28,
    2764 => -28,
    2765 => -28,
    2766 => -28,
    2767 => -28,
    2768 => -28,
    2769 => -28,
    2770 => -28,
    2771 => -28,
    2772 => -28,
    2773 => -28,
    2774 => -28,
    2775 => -28,
    2776 => -28,
    2777 => -28,
    2778 => -28,
    2779 => -28,
    2780 => -28,
    2781 => -28,
    2782 => -28,
    2783 => -29,
    2784 => -29,
    2785 => -29,
    2786 => -29,
    2787 => -29,
    2788 => -29,
    2789 => -29,
    2790 => -29,
    2791 => -29,
    2792 => -29,
    2793 => -29,
    2794 => -29,
    2795 => -29,
    2796 => -29,
    2797 => -29,
    2798 => -29,
    2799 => -29,
    2800 => -29,
    2801 => -29,
    2802 => -29,
    2803 => -29,
    2804 => -29,
    2805 => -29,
    2806 => -29,
    2807 => -29,
    2808 => -29,
    2809 => -29,
    2810 => -29,
    2811 => -29,
    2812 => -29,
    2813 => -29,
    2814 => -29,
    2815 => -29,
    2816 => -29,
    2817 => -29,
    2818 => -29,
    2819 => -29,
    2820 => -29,
    2821 => -29,
    2822 => -29,
    2823 => -29,
    2824 => -29,
    2825 => -29,
    2826 => -29,
    2827 => -29,
    2828 => -29,
    2829 => -29,
    2830 => -29,
    2831 => -29,
    2832 => -29,
    2833 => -29,
    2834 => -29,
    2835 => -29,
    2836 => -29,
    2837 => -30,
    2838 => -30,
    2839 => -30,
    2840 => -30,
    2841 => -30,
    2842 => -30,
    2843 => -30,
    2844 => -30,
    2845 => -30,
    2846 => -30,
    2847 => -30,
    2848 => -30,
    2849 => -30,
    2850 => -30,
    2851 => -30,
    2852 => -30,
    2853 => -30,
    2854 => -30,
    2855 => -30,
    2856 => -30,
    2857 => -30,
    2858 => -30,
    2859 => -30,
    2860 => -30,
    2861 => -30,
    2862 => -30,
    2863 => -30,
    2864 => -30,
    2865 => -30,
    2866 => -30,
    2867 => -30,
    2868 => -30,
    2869 => -30,
    2870 => -30,
    2871 => -30,
    2872 => -30,
    2873 => -30,
    2874 => -30,
    2875 => -30,
    2876 => -30,
    2877 => -30,
    2878 => -30,
    2879 => -30,
    2880 => -30,
    2881 => -30,
    2882 => -30,
    2883 => -30,
    2884 => -30,
    2885 => -30,
    2886 => -30,
    2887 => -30,
    2888 => -30,
    2889 => -30,
    2890 => -30,
    2891 => -30,
    2892 => -30,
    2893 => -30,
    2894 => -30,
    2895 => -30,
    2896 => -30,
    2897 => -30,
    2898 => -30,
    2899 => -30,
    2900 => -30,
    2901 => -30,
    2902 => -30,
    2903 => -30,
    2904 => -30,
    2905 => -30,
    2906 => -31,
    2907 => -31,
    2908 => -31,
    2909 => -31,
    2910 => -31,
    2911 => -31,
    2912 => -31,
    2913 => -31,
    2914 => -31,
    2915 => -31,
    2916 => -31,
    2917 => -31,
    2918 => -31,
    2919 => -31,
    2920 => -31,
    2921 => -31,
    2922 => -31,
    2923 => -31,
    2924 => -31,
    2925 => -31,
    2926 => -31,
    2927 => -31,
    2928 => -31,
    2929 => -31,
    2930 => -31,
    2931 => -31,
    2932 => -31,
    2933 => -31,
    2934 => -31,
    2935 => -31,
    2936 => -31,
    2937 => -31,
    2938 => -31,
    2939 => -31,
    2940 => -31,
    2941 => -31,
    2942 => -31,
    2943 => -31,
    2944 => -31,
    2945 => -31,
    2946 => -31,
    2947 => -31,
    2948 => -31,
    2949 => -31,
    2950 => -31,
    2951 => -31,
    2952 => -31,
    2953 => -31,
    2954 => -31,
    2955 => -31,
    2956 => -31,
    2957 => -31,
    2958 => -31,
    2959 => -31,
    2960 => -31,
    2961 => -31,
    2962 => -31,
    2963 => -31,
    2964 => -31,
    2965 => -31,
    2966 => -31,
    2967 => -31,
    2968 => -31,
    2969 => -31,
    2970 => -31,
    2971 => -31,
    2972 => -31,
    2973 => -31,
    2974 => -31,
    2975 => -31,
    2976 => -31,
    2977 => -31,
    2978 => -31,
    2979 => -31,
    2980 => -31,
    2981 => -31,
    2982 => -31,
    2983 => -31,
    2984 => -31,
    2985 => -31,
    2986 => -31,
    2987 => -31,
    2988 => -31,
    2989 => -31,
    2990 => -31,
    2991 => -31,
    2992 => -31,
    2993 => -31,
    2994 => -31,
    2995 => -31,
    2996 => -31,
    2997 => -31,
    2998 => -31,
    2999 => -31,
    3000 => -31,
    3001 => -31,
    3002 => -31,
    3003 => -31,
    3004 => -31,
    3005 => -31,
    3006 => -31,
    3007 => -31,
    3008 => -31,
    3009 => -31,
    3010 => -31,
    3011 => -31,
    3012 => -31,
    3013 => -31,
    3014 => -31,
    3015 => -31,
    3016 => -31,
    3017 => -31,
    3018 => -31,
    3019 => -31,
    3020 => -31,
    3021 => -31,
    3022 => -31,
    3023 => -31,
    3024 => -31,
    3025 => -31,
    3026 => -31,
    3027 => -31,
    3028 => -31,
    3029 => -31,
    3030 => -31,
    3031 => -31,
    3032 => -31,
    3033 => -31,
    3034 => -31,
    3035 => -31,
    3036 => -31,
    3037 => -31,
    3038 => -31,
    3039 => -31,
    3040 => -31,
    3041 => -31,
    3042 => -31,
    3043 => -31,
    3044 => -31,
    3045 => -31,
    3046 => -31,
    3047 => -31,
    3048 => -31,
    3049 => -31,
    3050 => -31,
    3051 => -31,
    3052 => -31,
    3053 => -31,
    3054 => -31,
    3055 => -31,
    3056 => -31,
    3057 => -31,
    3058 => -31,
    3059 => -31,
    3060 => -31,
    3061 => -31,
    3062 => -31,
    3063 => -31,
    3064 => -31,
    3065 => -31,
    3066 => -31,
    3067 => -31,
    3068 => -31,
    3069 => -31,
    3070 => -31,
    3071 => -31,
    3072 => -31,
    3073 => -31,
    3074 => -31,
    3075 => -31,
    3076 => -31,
    3077 => -31,
    3078 => -31,
    3079 => -31,
    3080 => -31,
    3081 => -31,
    3082 => -31,
    3083 => -31,
    3084 => -31,
    3085 => -31,
    3086 => -31,
    3087 => -31,
    3088 => -31,
    3089 => -31,
    3090 => -31,
    3091 => -31,
    3092 => -31,
    3093 => -31,
    3094 => -31,
    3095 => -31,
    3096 => -31,
    3097 => -31,
    3098 => -31,
    3099 => -31,
    3100 => -31,
    3101 => -31,
    3102 => -31,
    3103 => -31,
    3104 => -31,
    3105 => -31,
    3106 => -31,
    3107 => -31,
    3108 => -31,
    3109 => -31,
    3110 => -31,
    3111 => -31,
    3112 => -31,
    3113 => -31,
    3114 => -31,
    3115 => -31,
    3116 => -31,
    3117 => -31,
    3118 => -31,
    3119 => -31,
    3120 => -31,
    3121 => -31,
    3122 => -31,
    3123 => -31,
    3124 => -31,
    3125 => -31,
    3126 => -31,
    3127 => -31,
    3128 => -31,
    3129 => -31,
    3130 => -31,
    3131 => -31,
    3132 => -31,
    3133 => -31,
    3134 => -31,
    3135 => -31,
    3136 => -31,
    3137 => -31,
    3138 => -31,
    3139 => -31,
    3140 => -31,
    3141 => -31,
    3142 => -31,
    3143 => -31,
    3144 => -31,
    3145 => -31,
    3146 => -31,
    3147 => -31,
    3148 => -31,
    3149 => -31,
    3150 => -31,
    3151 => -31,
    3152 => -31,
    3153 => -31,
    3154 => -31,
    3155 => -31,
    3156 => -31,
    3157 => -31,
    3158 => -31,
    3159 => -31,
    3160 => -31,
    3161 => -31,
    3162 => -31,
    3163 => -31,
    3164 => -31,
    3165 => -31,
    3166 => -31,
    3167 => -31,
    3168 => -31,
    3169 => -31,
    3170 => -31,
    3171 => -31,
    3172 => -31,
    3173 => -31,
    3174 => -31,
    3175 => -31,
    3176 => -31,
    3177 => -31,
    3178 => -31,
    3179 => -31,
    3180 => -31,
    3181 => -31,
    3182 => -31,
    3183 => -31,
    3184 => -31,
    3185 => -31,
    3186 => -31,
    3187 => -31,
    3188 => -31,
    3189 => -31,
    3190 => -31,
    3191 => -31,
    3192 => -31,
    3193 => -31,
    3194 => -31,
    3195 => -31,
    3196 => -31,
    3197 => -31,
    3198 => -31,
    3199 => -31,
    3200 => -31,
    3201 => -31,
    3202 => -31,
    3203 => -31,
    3204 => -31,
    3205 => -31,
    3206 => -31,
    3207 => -31,
    3208 => -31,
    3209 => -31,
    3210 => -31,
    3211 => -31,
    3212 => -31,
    3213 => -31,
    3214 => -31,
    3215 => -31,
    3216 => -31,
    3217 => -31,
    3218 => -31,
    3219 => -31,
    3220 => -31,
    3221 => -31,
    3222 => -31,
    3223 => -31,
    3224 => -31,
    3225 => -31,
    3226 => -31,
    3227 => -31,
    3228 => -31,
    3229 => -31,
    3230 => -31,
    3231 => -31,
    3232 => -31,
    3233 => -31,
    3234 => -31,
    3235 => -31,
    3236 => -31,
    3237 => -31,
    3238 => -31,
    3239 => -30,
    3240 => -30,
    3241 => -30,
    3242 => -30,
    3243 => -30,
    3244 => -30,
    3245 => -30,
    3246 => -30,
    3247 => -30,
    3248 => -30,
    3249 => -30,
    3250 => -30,
    3251 => -30,
    3252 => -30,
    3253 => -30,
    3254 => -30,
    3255 => -30,
    3256 => -30,
    3257 => -30,
    3258 => -30,
    3259 => -30,
    3260 => -30,
    3261 => -30,
    3262 => -30,
    3263 => -30,
    3264 => -30,
    3265 => -30,
    3266 => -30,
    3267 => -30,
    3268 => -30,
    3269 => -30,
    3270 => -30,
    3271 => -30,
    3272 => -30,
    3273 => -30,
    3274 => -30,
    3275 => -30,
    3276 => -30,
    3277 => -30,
    3278 => -30,
    3279 => -30,
    3280 => -30,
    3281 => -30,
    3282 => -30,
    3283 => -30,
    3284 => -30,
    3285 => -30,
    3286 => -30,
    3287 => -30,
    3288 => -30,
    3289 => -30,
    3290 => -30,
    3291 => -30,
    3292 => -30,
    3293 => -30,
    3294 => -30,
    3295 => -30,
    3296 => -30,
    3297 => -30,
    3298 => -30,
    3299 => -30,
    3300 => -30,
    3301 => -30,
    3302 => -30,
    3303 => -30,
    3304 => -30,
    3305 => -30,
    3306 => -30,
    3307 => -30,
    3308 => -29,
    3309 => -29,
    3310 => -29,
    3311 => -29,
    3312 => -29,
    3313 => -29,
    3314 => -29,
    3315 => -29,
    3316 => -29,
    3317 => -29,
    3318 => -29,
    3319 => -29,
    3320 => -29,
    3321 => -29,
    3322 => -29,
    3323 => -29,
    3324 => -29,
    3325 => -29,
    3326 => -29,
    3327 => -29,
    3328 => -29,
    3329 => -29,
    3330 => -29,
    3331 => -29,
    3332 => -29,
    3333 => -29,
    3334 => -29,
    3335 => -29,
    3336 => -29,
    3337 => -29,
    3338 => -29,
    3339 => -29,
    3340 => -29,
    3341 => -29,
    3342 => -29,
    3343 => -29,
    3344 => -29,
    3345 => -29,
    3346 => -29,
    3347 => -29,
    3348 => -29,
    3349 => -29,
    3350 => -29,
    3351 => -29,
    3352 => -29,
    3353 => -29,
    3354 => -29,
    3355 => -29,
    3356 => -29,
    3357 => -29,
    3358 => -29,
    3359 => -29,
    3360 => -29,
    3361 => -29,
    3362 => -28,
    3363 => -28,
    3364 => -28,
    3365 => -28,
    3366 => -28,
    3367 => -28,
    3368 => -28,
    3369 => -28,
    3370 => -28,
    3371 => -28,
    3372 => -28,
    3373 => -28,
    3374 => -28,
    3375 => -28,
    3376 => -28,
    3377 => -28,
    3378 => -28,
    3379 => -28,
    3380 => -28,
    3381 => -28,
    3382 => -28,
    3383 => -28,
    3384 => -28,
    3385 => -28,
    3386 => -28,
    3387 => -28,
    3388 => -28,
    3389 => -28,
    3390 => -28,
    3391 => -28,
    3392 => -28,
    3393 => -28,
    3394 => -28,
    3395 => -28,
    3396 => -28,
    3397 => -28,
    3398 => -28,
    3399 => -28,
    3400 => -28,
    3401 => -28,
    3402 => -28,
    3403 => -28,
    3404 => -28,
    3405 => -28,
    3406 => -28,
    3407 => -27,
    3408 => -27,
    3409 => -27,
    3410 => -27,
    3411 => -27,
    3412 => -27,
    3413 => -27,
    3414 => -27,
    3415 => -27,
    3416 => -27,
    3417 => -27,
    3418 => -27,
    3419 => -27,
    3420 => -27,
    3421 => -27,
    3422 => -27,
    3423 => -27,
    3424 => -27,
    3425 => -27,
    3426 => -27,
    3427 => -27,
    3428 => -27,
    3429 => -27,
    3430 => -27,
    3431 => -27,
    3432 => -27,
    3433 => -27,
    3434 => -27,
    3435 => -27,
    3436 => -27,
    3437 => -27,
    3438 => -27,
    3439 => -27,
    3440 => -27,
    3441 => -27,
    3442 => -27,
    3443 => -27,
    3444 => -27,
    3445 => -27,
    3446 => -27,
    3447 => -27,
    3448 => -26,
    3449 => -26,
    3450 => -26,
    3451 => -26,
    3452 => -26,
    3453 => -26,
    3454 => -26,
    3455 => -26,
    3456 => -26,
    3457 => -26,
    3458 => -26,
    3459 => -26,
    3460 => -26,
    3461 => -26,
    3462 => -26,
    3463 => -26,
    3464 => -26,
    3465 => -26,
    3466 => -26,
    3467 => -26,
    3468 => -26,
    3469 => -26,
    3470 => -26,
    3471 => -26,
    3472 => -26,
    3473 => -26,
    3474 => -26,
    3475 => -26,
    3476 => -26,
    3477 => -26,
    3478 => -26,
    3479 => -26,
    3480 => -26,
    3481 => -26,
    3482 => -26,
    3483 => -26,
    3484 => -26,
    3485 => -25,
    3486 => -25,
    3487 => -25,
    3488 => -25,
    3489 => -25,
    3490 => -25,
    3491 => -25,
    3492 => -25,
    3493 => -25,
    3494 => -25,
    3495 => -25,
    3496 => -25,
    3497 => -25,
    3498 => -25,
    3499 => -25,
    3500 => -25,
    3501 => -25,
    3502 => -25,
    3503 => -25,
    3504 => -25,
    3505 => -25,
    3506 => -25,
    3507 => -25,
    3508 => -25,
    3509 => -25,
    3510 => -25,
    3511 => -25,
    3512 => -25,
    3513 => -25,
    3514 => -25,
    3515 => -25,
    3516 => -25,
    3517 => -25,
    3518 => -25,
    3519 => -24,
    3520 => -24,
    3521 => -24,
    3522 => -24,
    3523 => -24,
    3524 => -24,
    3525 => -24,
    3526 => -24,
    3527 => -24,
    3528 => -24,
    3529 => -24,
    3530 => -24,
    3531 => -24,
    3532 => -24,
    3533 => -24,
    3534 => -24,
    3535 => -24,
    3536 => -24,
    3537 => -24,
    3538 => -24,
    3539 => -24,
    3540 => -24,
    3541 => -24,
    3542 => -24,
    3543 => -24,
    3544 => -24,
    3545 => -24,
    3546 => -24,
    3547 => -24,
    3548 => -24,
    3549 => -24,
    3550 => -24,
    3551 => -24,
    3552 => -23,
    3553 => -23,
    3554 => -23,
    3555 => -23,
    3556 => -23,
    3557 => -23,
    3558 => -23,
    3559 => -23,
    3560 => -23,
    3561 => -23,
    3562 => -23,
    3563 => -23,
    3564 => -23,
    3565 => -23,
    3566 => -23,
    3567 => -23,
    3568 => -23,
    3569 => -23,
    3570 => -23,
    3571 => -23,
    3572 => -23,
    3573 => -23,
    3574 => -23,
    3575 => -23,
    3576 => -23,
    3577 => -23,
    3578 => -23,
    3579 => -23,
    3580 => -23,
    3581 => -23,
    3582 => -22,
    3583 => -22,
    3584 => -22,
    3585 => -22,
    3586 => -22,
    3587 => -22,
    3588 => -22,
    3589 => -22,
    3590 => -22,
    3591 => -22,
    3592 => -22,
    3593 => -22,
    3594 => -22,
    3595 => -22,
    3596 => -22,
    3597 => -22,
    3598 => -22,
    3599 => -22,
    3600 => -22,
    3601 => -22,
    3602 => -22,
    3603 => -22,
    3604 => -22,
    3605 => -22,
    3606 => -22,
    3607 => -22,
    3608 => -22,
    3609 => -22,
    3610 => -22,
    3611 => -21,
    3612 => -21,
    3613 => -21,
    3614 => -21,
    3615 => -21,
    3616 => -21,
    3617 => -21,
    3618 => -21,
    3619 => -21,
    3620 => -21,
    3621 => -21,
    3622 => -21,
    3623 => -21,
    3624 => -21,
    3625 => -21,
    3626 => -21,
    3627 => -21,
    3628 => -21,
    3629 => -21,
    3630 => -21,
    3631 => -21,
    3632 => -21,
    3633 => -21,
    3634 => -21,
    3635 => -21,
    3636 => -21,
    3637 => -21,
    3638 => -21,
    3639 => -20,
    3640 => -20,
    3641 => -20,
    3642 => -20,
    3643 => -20,
    3644 => -20,
    3645 => -20,
    3646 => -20,
    3647 => -20,
    3648 => -20,
    3649 => -20,
    3650 => -20,
    3651 => -20,
    3652 => -20,
    3653 => -20,
    3654 => -20,
    3655 => -20,
    3656 => -20,
    3657 => -20,
    3658 => -20,
    3659 => -20,
    3660 => -20,
    3661 => -20,
    3662 => -20,
    3663 => -20,
    3664 => -20,
    3665 => -20,
    3666 => -19,
    3667 => -19,
    3668 => -19,
    3669 => -19,
    3670 => -19,
    3671 => -19,
    3672 => -19,
    3673 => -19,
    3674 => -19,
    3675 => -19,
    3676 => -19,
    3677 => -19,
    3678 => -19,
    3679 => -19,
    3680 => -19,
    3681 => -19,
    3682 => -19,
    3683 => -19,
    3684 => -19,
    3685 => -19,
    3686 => -19,
    3687 => -19,
    3688 => -19,
    3689 => -19,
    3690 => -19,
    3691 => -19,
    3692 => -19,
    3693 => -18,
    3694 => -18,
    3695 => -18,
    3696 => -18,
    3697 => -18,
    3698 => -18,
    3699 => -18,
    3700 => -18,
    3701 => -18,
    3702 => -18,
    3703 => -18,
    3704 => -18,
    3705 => -18,
    3706 => -18,
    3707 => -18,
    3708 => -18,
    3709 => -18,
    3710 => -18,
    3711 => -18,
    3712 => -18,
    3713 => -18,
    3714 => -18,
    3715 => -18,
    3716 => -18,
    3717 => -18,
    3718 => -17,
    3719 => -17,
    3720 => -17,
    3721 => -17,
    3722 => -17,
    3723 => -17,
    3724 => -17,
    3725 => -17,
    3726 => -17,
    3727 => -17,
    3728 => -17,
    3729 => -17,
    3730 => -17,
    3731 => -17,
    3732 => -17,
    3733 => -17,
    3734 => -17,
    3735 => -17,
    3736 => -17,
    3737 => -17,
    3738 => -17,
    3739 => -17,
    3740 => -17,
    3741 => -17,
    3742 => -17,
    3743 => -16,
    3744 => -16,
    3745 => -16,
    3746 => -16,
    3747 => -16,
    3748 => -16,
    3749 => -16,
    3750 => -16,
    3751 => -16,
    3752 => -16,
    3753 => -16,
    3754 => -16,
    3755 => -16,
    3756 => -16,
    3757 => -16,
    3758 => -16,
    3759 => -16,
    3760 => -16,
    3761 => -16,
    3762 => -16,
    3763 => -16,
    3764 => -16,
    3765 => -16,
    3766 => -16,
    3767 => -15,
    3768 => -15,
    3769 => -15,
    3770 => -15,
    3771 => -15,
    3772 => -15,
    3773 => -15,
    3774 => -15,
    3775 => -15,
    3776 => -15,
    3777 => -15,
    3778 => -15,
    3779 => -15,
    3780 => -15,
    3781 => -15,
    3782 => -15,
    3783 => -15,
    3784 => -15,
    3785 => -15,
    3786 => -15,
    3787 => -15,
    3788 => -15,
    3789 => -15,
    3790 => -15,
    3791 => -14,
    3792 => -14,
    3793 => -14,
    3794 => -14,
    3795 => -14,
    3796 => -14,
    3797 => -14,
    3798 => -14,
    3799 => -14,
    3800 => -14,
    3801 => -14,
    3802 => -14,
    3803 => -14,
    3804 => -14,
    3805 => -14,
    3806 => -14,
    3807 => -14,
    3808 => -14,
    3809 => -14,
    3810 => -14,
    3811 => -14,
    3812 => -14,
    3813 => -14,
    3814 => -13,
    3815 => -13,
    3816 => -13,
    3817 => -13,
    3818 => -13,
    3819 => -13,
    3820 => -13,
    3821 => -13,
    3822 => -13,
    3823 => -13,
    3824 => -13,
    3825 => -13,
    3826 => -13,
    3827 => -13,
    3828 => -13,
    3829 => -13,
    3830 => -13,
    3831 => -13,
    3832 => -13,
    3833 => -13,
    3834 => -13,
    3835 => -13,
    3836 => -13,
    3837 => -12,
    3838 => -12,
    3839 => -12,
    3840 => -12,
    3841 => -12,
    3842 => -12,
    3843 => -12,
    3844 => -12,
    3845 => -12,
    3846 => -12,
    3847 => -12,
    3848 => -12,
    3849 => -12,
    3850 => -12,
    3851 => -12,
    3852 => -12,
    3853 => -12,
    3854 => -12,
    3855 => -12,
    3856 => -12,
    3857 => -12,
    3858 => -12,
    3859 => -12,
    3860 => -11,
    3861 => -11,
    3862 => -11,
    3863 => -11,
    3864 => -11,
    3865 => -11,
    3866 => -11,
    3867 => -11,
    3868 => -11,
    3869 => -11,
    3870 => -11,
    3871 => -11,
    3872 => -11,
    3873 => -11,
    3874 => -11,
    3875 => -11,
    3876 => -11,
    3877 => -11,
    3878 => -11,
    3879 => -11,
    3880 => -11,
    3881 => -11,
    3882 => -10,
    3883 => -10,
    3884 => -10,
    3885 => -10,
    3886 => -10,
    3887 => -10,
    3888 => -10,
    3889 => -10,
    3890 => -10,
    3891 => -10,
    3892 => -10,
    3893 => -10,
    3894 => -10,
    3895 => -10,
    3896 => -10,
    3897 => -10,
    3898 => -10,
    3899 => -10,
    3900 => -10,
    3901 => -10,
    3902 => -10,
    3903 => -10,
    3904 => -9,
    3905 => -9,
    3906 => -9,
    3907 => -9,
    3908 => -9,
    3909 => -9,
    3910 => -9,
    3911 => -9,
    3912 => -9,
    3913 => -9,
    3914 => -9,
    3915 => -9,
    3916 => -9,
    3917 => -9,
    3918 => -9,
    3919 => -9,
    3920 => -9,
    3921 => -9,
    3922 => -9,
    3923 => -9,
    3924 => -9,
    3925 => -9,
    3926 => -8,
    3927 => -8,
    3928 => -8,
    3929 => -8,
    3930 => -8,
    3931 => -8,
    3932 => -8,
    3933 => -8,
    3934 => -8,
    3935 => -8,
    3936 => -8,
    3937 => -8,
    3938 => -8,
    3939 => -8,
    3940 => -8,
    3941 => -8,
    3942 => -8,
    3943 => -8,
    3944 => -8,
    3945 => -8,
    3946 => -8,
    3947 => -8,
    3948 => -7,
    3949 => -7,
    3950 => -7,
    3951 => -7,
    3952 => -7,
    3953 => -7,
    3954 => -7,
    3955 => -7,
    3956 => -7,
    3957 => -7,
    3958 => -7,
    3959 => -7,
    3960 => -7,
    3961 => -7,
    3962 => -7,
    3963 => -7,
    3964 => -7,
    3965 => -7,
    3966 => -7,
    3967 => -7,
    3968 => -7,
    3969 => -7,
    3970 => -6,
    3971 => -6,
    3972 => -6,
    3973 => -6,
    3974 => -6,
    3975 => -6,
    3976 => -6,
    3977 => -6,
    3978 => -6,
    3979 => -6,
    3980 => -6,
    3981 => -6,
    3982 => -6,
    3983 => -6,
    3984 => -6,
    3985 => -6,
    3986 => -6,
    3987 => -6,
    3988 => -6,
    3989 => -6,
    3990 => -6,
    3991 => -5,
    3992 => -5,
    3993 => -5,
    3994 => -5,
    3995 => -5,
    3996 => -5,
    3997 => -5,
    3998 => -5,
    3999 => -5,
    4000 => -5,
    4001 => -5,
    4002 => -5,
    4003 => -5,
    4004 => -5,
    4005 => -5,
    4006 => -5,
    4007 => -5,
    4008 => -5,
    4009 => -5,
    4010 => -5,
    4011 => -5,
    4012 => -4,
    4013 => -4,
    4014 => -4,
    4015 => -4,
    4016 => -4,
    4017 => -4,
    4018 => -4,
    4019 => -4,
    4020 => -4,
    4021 => -4,
    4022 => -4,
    4023 => -4,
    4024 => -4,
    4025 => -4,
    4026 => -4,
    4027 => -4,
    4028 => -4,
    4029 => -4,
    4030 => -4,
    4031 => -4,
    4032 => -4,
    4033 => -3,
    4034 => -3,
    4035 => -3,
    4036 => -3,
    4037 => -3,
    4038 => -3,
    4039 => -3,
    4040 => -3,
    4041 => -3,
    4042 => -3,
    4043 => -3,
    4044 => -3,
    4045 => -3,
    4046 => -3,
    4047 => -3,
    4048 => -3,
    4049 => -3,
    4050 => -3,
    4051 => -3,
    4052 => -3,
    4053 => -3,
    4054 => -2,
    4055 => -2,
    4056 => -2,
    4057 => -2,
    4058 => -2,
    4059 => -2,
    4060 => -2,
    4061 => -2,
    4062 => -2,
    4063 => -2,
    4064 => -2,
    4065 => -2,
    4066 => -2,
    4067 => -2,
    4068 => -2,
    4069 => -2,
    4070 => -2,
    4071 => -2,
    4072 => -2,
    4073 => -2,
    4074 => -2,
    4075 => -1,
    4076 => -1,
    4077 => -1,
    4078 => -1,
    4079 => -1,
    4080 => -1,
    4081 => -1,
    4082 => -1,
    4083 => -1,
    4084 => -1,
    4085 => -1,
    4086 => -1,
    4087 => -1,
    4088 => -1,
    4089 => -1,
    4090 => -1,
    4091 => -1,
    4092 => -1,
    4093 => -1,
    4094 => -1,
    4095 => -1
);

begin
  dds_out <= std_logic_vector(TO_SIGNED(LUT(TO_INTEGER(unsigned(address))),6));
end rtl;
