library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all; -- for the casting 
	
-- This testbench aims to check if the output
-- of the filter is the same as the one designed in MATLAB

entity IIR_TB_Street is
end IIR_TB_Street;

architecture TB_Arch of IIR_TB_Street is	

component IIR  
	generic (Nbit : natural := 8);
	port (
		clk		:	in	std_logic;
		rst_l	:	in	std_logic;
		x		:	in	std_logic_vector(Nbit-1 downto 0);	
		y		:	out	std_logic_vector(Nbit-1 downto 0)
	);
end component;

	constant BITS		:	natural	:=	16;
	constant SAMPLES 	:	natural	:= 	1000;

	signal clk		: 	std_logic	:= '0'; -- initial value. It's not something physically possible to initialize it but in testbench is ok 
	signal rst_l 	: 	std_logic;
	signal sample	:	std_logic_vector(BITS-1 downto 0);
	signal output	:	std_logic_vector(BITS-1 downto 0);
	signal expected	:	std_logic_vector(BITS-1 downto 0);
	
	signal enable	:	std_logic	:=	'1';
	
	-- Data type to store the sequence of samples
	type WAV_IN is array (0 to SAMPLES-1) of std_logic_vector(BITS-1 downto 0);

begin
	
	filter: IIR
	generic map(BITS)
	port map(clk, rst_l, sample, output);
	
	-- clock generator
	clk <= not clk and enable after 11338 ns; -- 44100Hz clock
	
	-- stimuli
	driver_p: process
	
	variable input : WAV_IN := ("1111111111100011",
								"0000000001001100",
								"0000000011111110",
								"0000000100011001",
								"0000000011101101",
								"0000000100111001",
								"0000000011101111",
								"0000000011110100",
								"0000000100000010",
								"0000000011000110",
								"0000000000001000",
								"1111111111010101",
								"1111111111111010",
								"1111111111001101",
								"0000000010010100",
								"0000000011000010",
								"0000000110001100",
								"0000000111111100",
								"0000001001000000",
								"0000001001010010",
								"0000001010111110",
								"0000001101011001",
								"0000001100110110",
								"0000001110100000",
								"0000001110110100",
								"0000001111111101",
								"0000010000011110",
								"0000010001100000",
								"0000010010010001",
								"0000010011001001",
								"0000010011010010",
								"0000010100011011",
								"0000010100110100",
								"0000010101101000",
								"0000010100110010",
								"0000010101100010",
								"0000010111111110",
								"0000010111101011",
								"0000011000001011",
								"0000011001001100",
								"0000011001101101",
								"0000011010001110",
								"0000011010010010",
								"0000011011100110",
								"0000011011101101",
								"0000011101011110",
								"0000100000110111",
								"0000100010101000",
								"0000100001100111",
								"0000100011011011",
								"0000100011010100",
								"0000100100000011",
								"0000100011101101",
								"0000100100000111",
								"0000100010001010",
								"0000100000111111",
								"0000100001110011",
								"0000100010010000",
								"0000100011011011",
								"0000100011101000",
								"0000100011010111",
								"0000100100000111",
								"0000100100010000",
								"0000100100001010",
								"0000100100010100",
								"0000100101111110",
								"0000100101011111",
								"0000100101111111",
								"0000100110010100",
								"0000100111001011",
								"0000100110111001",
								"0000100111111110",
								"0000100111110011",
								"0000101000101100",
								"0000101000100101",
								"0000101000111000",
								"0000100110101110",
								"0000100011011100",
								"0000100101000111",
								"0000100101101001",
								"0000100101011100",
								"0000100110001001",
								"0000100101111101",
								"0000100110101100",
								"0000100110000000",
								"0000100110010101",
								"0000100110000001",
								"0000100110011000",
								"0000100110010111",
								"0000100111100110",
								"0000101010001100",
								"0000101011000011",
								"0000101010000111",
								"0000101010110111",
								"0000101001110010",
								"0000101010001111",
								"0000101001101001",
								"0000101001001010",
								"0000100110110010",
								"0000100101010111",
								"0000100100001101",
								"0000100100110011",
								"0000100100100101",
								"0000100011101010",
								"0000100100101111",
								"0000100011011010",
								"0000100011111111",
								"0000100010001111",
								"0000100011000101",
								"0000100011001100",
								"0000100010011000",
								"0000100010101100",
								"0000100010001011",
								"0000100010001011",
								"0000100001110001",
								"0000100001111010",
								"0000100001101110",
								"0000100010101111",
								"0000110110101010",
								"0001011011000010",
								"0001010000101010",
								"0001000101010010",
								"0001001011100010",
								"0000111111110011",
								"0001000101101101",
								"0000111101111011",
								"0001000001010011",
								"0000111100110011",
								"0000111110110100",
								"0000111100000000",
								"0000111101011000",
								"0000111011101100",
								"0000111100101000",
								"0000111100001101",
								"0000111111110011",
								"0001000000110001",
								"0001000000000010",
								"0001000000100010",
								"0001000000100011",
								"0001000000011111",
								"0000111111111010",
								"0001000000000100",
								"0000111101110110",
								"0000111100000101",
								"0000111011111010",
								"0000111011110110",
								"0000111100100000",
								"0000111100111100",
								"0000111100011011",
								"0000111100111101",
								"0000111100111010",
								"0000111100100000",
								"0000111100010100",
								"0000111101110101",
								"0000111100101001",
								"0000111101010101",
								"0000111101001001",
								"0000111110000001",
								"0000111100101000",
								"0000100101001010",
								"1110110100001000",
								"1110000111110110",
								"1111100101001001",
								"1111010100011000",
								"1111110000101001",
								"1111111000001000",
								"1111111001100110",
								"0000000111011000",
								"0000000000000101",
								"0000001110000000",
								"0000000100000001",
								"0000010000111000",
								"0000000111001100",
								"0000010010100110",
								"0000001000101010",
								"0000010010110001",
								"0000001010100001",
								"0000010011101110",
								"0000001110111011",
								"0000011000001100",
								"0000010000010011",
								"0000010111101010",
								"0000010010000000",
								"0000010110111101",
								"0000010010000011",
								"0000010110010011",
								"0000010000011101",
								"0000010010001111",
								"0000001111000010",
								"0000010010010001",
								"0000001110101011",
								"0000010010010110",
								"0000001111000101",
								"0000010010111110",
								"0000001111011010",
								"0000010001010110",
								"0000001110111101",
								"0000010010100011",
								"0000001111001010",
								"0000010001110001",
								"0000001111011001",
								"0000011101110111",
								"0001111001011110",
								"0011011011000100",
								"0010010010011010",
								"0010001101101010",
								"0010001000111111",
								"0001101111100101",
								"0001111001010111",
								"0001100001110010",
								"0001101100011010",
								"0001011010001010",
								"0001100011001111",
								"0001010101010001",
								"0001011100111011",
								"0001010010110101",
								"0001010111111000",
								"0001010001000011",
								"0001010100100101",
								"0001001111011110",
								"0001010010001111",
								"0001001110110010",
								"0001010011111110",
								"0001010011010001",
								"0001010011100110",
								"0001010001011110",
								"0001010011011101",
								"0001010000010011",
								"0001010010010010",
								"0001010000000001",
								"0001001111011011",
								"0001001011001111",
								"0001001100110000",
								"0001001011001110",
								"0001001011111010",
								"0001001010100010",
								"0001001011101000",
								"0001001010100111",
								"0001001011011111",
								"0001001001011001",
								"0001001001110100",
								"0001001010100101",
								"0001000111101110",
								"1111110010100111",
								"1011110111100101",
								"1011111011011111",
								"1110101000001100",
								"1101110001111111",
								"1111001011011101",
								"1110110111001001",
								"1111011010010000",
								"1111011001111100",
								"1111100010100100",
								"1111101011110010",
								"1111101000000000",
								"1111110100010101",
								"1111101011111010",
								"1111111001011000",
								"1111101110101101",
								"1111111100001000",
								"1111110000010101",
								"1111111110001100",
								"1111110010100001",
								"1111111111000010",
								"1111110100000100",
								"1111111111111000",
								"1111111000100010",
								"0000000101111110",
								"1111111011010011",
								"0000000101101110",
								"1111111100111111",
								"0000000101110110",
								"1111111101101100",
								"0000000101110101",
								"1111111100110000",
								"0000000010010010",
								"1111111010010101",
								"0000000010110010",
								"1111111011111101",
								"0000000010111011",
								"1111111100010111",
								"0000000010110101",
								"1111111101010010",
								"0000000011000001",
								"1111111100110001",
								"0000100110111100",
								"0011001111111011",
								"0100111011000010",
								"0010110110011110",
								"0011010000101001",
								"0010101010010111",
								"0010011011110101",
								"0010010111110001",
								"0010000000010000",
								"0010001000000111",
								"0001110000111010",
								"0001111011001000",
								"0001101000001111",
								"0001110010011000",
								"0001100010010011",
								"0001101011011110",
								"0001011110011101",
								"0001100110001100",
								"0001011011100010",
								"0001100010100101",
								"0001011001011010",
								"0001011111101001",
								"0001010111110011",
								"0001011101001000",
								"0001010111010000",
								"0001011101100111",
								"0001011010110011",
								"0001011110001011",
								"0001011001000111",
								"0001011101001000",
								"0001010111111010",
								"0001011011101011",
								"0001010110110010",
								"0001011000110101",
								"0001010010001100",
								"0001010100100110",
								"0001010001101011",
								"0001010100000011",
								"0001010001010110",
								"0001010010110000",
								"0001010000111101",
								"0001001001111110",
								"1110101011101101",
								"1001111100101000",
								"1011101111010101",
								"1110000110000011",
								"1101001100110101",
								"1111000100001101",
								"1110010010110111",
								"1111011001100010",
								"1110111010011011",
								"1111100001110100",
								"1111010001101000",
								"1111100110000110",
								"1111011110110010",
								"1111100111111111",
								"1111100110110000",
								"1111101001110010",
								"1111101011011000",
								"1111101010111110",
								"1111101111001111",
								"1111101100000001",
								"1111110001101011",
								"1111101100111011",
								"1111110011101111",
								"1111101110001111",
								"1111110100101000",
								"1111101111110111",
								"1111110110000000",
								"1111110010100000",
								"1111111100000110",
								"1111110110011011",
								"1111111100010001",
								"1111110111011100",
								"1111111101000010",
								"1111110111100111",
								"1111111101110001",
								"1111110111100001",
								"1111111010000011",
								"1111110101011111",
								"1111111010001111",
								"1111110101111010",
								"1111111010001000",
								"1111111000001011",
								"0001000111010011",
								"0100111001010101",
								"0101100111100010",
								"0011001101000001",
								"0100000101001000",
								"0010110110010100",
								"0011000011001001",
								"0010100010101110",
								"0010011101000010",
								"0010010010100110",
								"0010000101111111",
								"0010000110001011",
								"0001110110111110",
								"0001111100101011",
								"0001101101100001",
								"0001110100111110",
								"0001100111010011",
								"0001101111000010",
								"0001100010011110",
								"0001101010010111",
								"0001011110110101",
								"0001100110100010",
								"0001011100000000",
								"0001100011010010",
								"0001011001100101",
								"0001100000100100",
								"0001010111101101",
								"0001011101110110",
								"0001010110001111",
								"0001011101100011",
								"0001011000111001",
								"0001011110101010",
								"0001010111100000",
								"0001011101010111",
								"0001010101011011",
								"0001011011101011",
								"0001010100101010",
								"0001011000111010",
								"0001001111011001",
								"0001010011100101",
								"0001001110110111",
								"0000111010001011",
								"1101010100011100",
								"1001010110001110",
								"1100101101010100",
								"1101101001011011",
								"1101011111110110",
								"1110111111100011",
								"1110010000111011",
								"1111011111101010",
								"1110110001000010",
								"1111101011000010",
								"1111000110100100",
								"1111101111000000",
								"1111010010101100",
								"1111110001101100",
								"1111011011100011",
								"1111110001110010",
								"1111100001111111",
								"1111110010011011",
								"1111100101110001",
								"1111110010111101",
								"1111101001011100",
								"1111110011010111",
								"1111101100011011",
								"1111110011101100",
								"1111101110011100",
								"1111110100010101",
								"1111110000001000",
								"1111110100110100",
								"1111110001111111",
								"1111110101010000",
								"1111110011010100",
								"1111110111101101",
								"1111111000111100",
								"1111111011110111",
								"1111111001001001",
								"1111111100110101",
								"1111111010011100",
								"1111111100110110",
								"1111111011001001",
								"1111111100010101",
								"1111111000101011",
								"1111111111010111",
								"0001110110011100",
								"0101111000011110",
								"0101001001001011",
								"0011011010011011",
								"0100001001110000",
								"0010110010000000",
								"0011010000011100",
								"0010011011110010",
								"0010101001011010",
								"0010001110001011",
								"0010010000100000",
								"0010000010011110",
								"0010000000100011",
								"0001111010101001",
								"0001110101000011",
								"0001110011101100",
								"0001101101010001",
								"0001101110111000",
								"0001100111110010",
								"0001101010101011",
								"0001100011010110",
								"0001100111001001",
								"0001100000000111",
								"0001100100010001",
								"0001011101000010",
								"0001100001111011",
								"0001011010101001",
								"0001011111010001",
								"0001011000100111",
								"0001011101100101",
								"0001010111000011",
								"0001011010111010",
								"0001010101011110",
								"0001011011001101",
								"0001011000001000",
								"0001011100101110",
								"0001010110111011",
								"0001011011000011",
								"0001010110000001",
								"0001011001001101",
								"0001010100100111",
								"0000100101011011",
								"1100000001101111",
								"1001011111110110",
								"1101100011001010",
								"1101001110000100",
								"1110000100011011",
								"1110110001010111",
								"1110100010100100",
								"1111011001111010",
								"1110111000111100",
								"1111101010101011",
								"1111000110101101",
								"1111110010100001",
								"1111010001101000",
								"1111110101001010",
								"1111011000111011",
								"1111110110100100",
								"1111011110001111",
								"1111110111000100",
								"1111100010100111",
								"1111110111011001",
								"1111100110001011",
								"1111111000000011",
								"1111101000001011",
								"1111111000010011",
								"1111101010011111",
								"1111111000110101",
								"1111101100111101",
								"1111111000101001",
								"1111101110011000",
								"1111111001101001",
								"1111101111100110",
								"1111111010000001",
								"1111110001011101",
								"1111111001111010",
								"1111110010001110",
								"1111111011011100",
								"1111110111110100",
								"1111111111111010",
								"1111111000111111",
								"0000000000000101",
								"1111111001110100",
								"0000010000010010",
								"0010110101011010",
								"0110100011100001",
								"0100100001100101",
								"0011110001000001",
								"0011111110100010",
								"0010110101011000",
								"0011010010000110",
								"0010011001101111",
								"0010110000000001",
								"0010001001101111",
								"0010011000010001",
								"0001111101111000",
								"0010000111010010",
								"0001110111001100",
								"0001111011011110",
								"0001110001000110",
								"0001110011001011",
								"0001101100100111",
								"0001101100101111",
								"0001101000100000",
								"0001101000000010",
								"0001100101101000",
								"0001100100000111",
								"0001100010110010",
								"0001100000110001",
								"0001100000011000",
								"0001011110000110",
								"0001011110100010",
								"0001011011110000",
								"0001011100010011",
								"0001011010000011",
								"0001011010011001",
								"0001010111110011",
								"0001011000111111",
								"0001010110000101",
								"0001010111001100",
								"0001010100110101",
								"0001010110100000",
								"0001010111011000",
								"0001011001110011",
								"0001010011101001",
								"1111111011010100",
								"1010110101000000",
								"1010010000000010",
								"1110000100101010",
								"1101000000000000",
								"1110101001100111",
								"1110011011011100",
								"1110111011111011",
								"1111001010010011",
								"1111001001000111",
								"1111100000100001",
								"1111010001001110",
								"1111101100000110",
								"1111010111111110",
								"1111110001000101",
								"1111011011000111",
								"1111110100111011",
								"1111011111101011",
								"1111110110010101",
								"1111100010011010",
								"1111110111100000",
								"1111100101011101",
								"1111111000001110",
								"1111100111110101",
								"1111111000110100",
								"1111101001101100",
								"1111111001001100",
								"1111101011100010",
								"1111111001100001",
								"1111101101001101",
								"1111111010001001",
								"1111101110001110",
								"1111111011000000",
								"1111101111100100",
								"1111111010110001",
								"1111110001000101",
								"1111111011001110",
								"1111110010000101",
								"1111111011100000",
								"1111110010111111",
								"1111111100100000",
								"1111110111000001",
								"0000100101100011",
								"0011111011000100",
								"0110101111010001",
								"0011111101100001",
								"0100001110000110",
								"0011101010010011",
								"0011000101111010",
								"0011001001001010",
								"0010011101001011",
								"0010101101000110",
								"0010001000100010",
								"0010011000111111",
								"0001111100011111",
								"0010001001111011",
								"0001110011101110",
								"0001111111101011",
								"0001101101011101",
								"0001110101111011",
								"0001101001010100",
								"0001110000000000",
								"0001100101010010",
								"0001101011010101",
								"0001100010000001",
								"0001100111010111",
								"0001011111010111",
								"0001100011110100",
								"0001011101011000",
								"0001100000100110",
								"0001011011011001",
								"0001011101110101",
								"0001011001110001",
								"0001011011100001",
								"0001010111110110",
								"0001011001011100",
								"0001010110011100",
								"0001010111101111",
								"0001010100101010",
								"0001010101101111",
								"0001010010111000",
								"0001010100100010",
								"0001010010011110",
								"0001001100101001",
								"1110111100110111",
								"1001110111110111",
								"1011001011100100",
								"1110000110111011",
								"1100111111011000",
								"1111000001011000",
								"1110010000100111",
								"1111010101010010",
								"1110111101011101",
								"1111011011010110",
								"1111010001101000",
								"1111011110001010",
								"1111011111100011",
								"1111100001101100",
								"1111100111100100",
								"1111100011001011",
								"1111101100101111",
								"1111100101101011",
								"1111101111100010",
								"1111100110000000",
								"1111110010110010",
								"1111101000101011",
								"1111110010100111",
								"1111101010101101",
								"1111110100000000",
								"1111101011011100",
								"1111110101011101",
								"1111101100100011",
								"1111110110001000",
								"1111101110001101",
								"1111110110100101",
								"1111101110101100",
								"1111110111111011",
								"1111101111111000",
								"1111111000000101",
								"1111110001001011",
								"1111111000010101",
								"1111110010001000",
								"1111111000110101",
								"1111110010110111",
								"1111111001000010",
								"1111110100011100",
								"0000110110100110",
								"0100110001011110",
								"0110011011000110",
								"0011101000100001",
								"0100011100001011",
								"0011010101001000",
								"0011010001001101",
								"0010111101111111",
								"0010101000000000",
								"0010101001011110",
								"0010001111010000",
								"0010010111010110",
								"0001111100100001",
								"0010000111111110",
								"0001110010010100",
								"0001111101100101",
								"0001101100000110",
								"0001110110001010",
								"0001100111011011",
								"0001110000101001",
								"0001100010111011",
								"0001101010011111",
								"0001011111111001",
								"0001100111101101",
								"0001011100101001",
								"0001100100011011",
								"0001011010010001",
								"0001100001001100",
								"0001011000100101",
								"0001011110010101",
								"0001010110011000",
								"0001011100000110",
								"0001010101001110",
								"0001011001011001",
								"0001010011011101",
								"0001010111100101",
								"0001010001100111",
								"0001010101111010",
								"0001010000101001",
								"0001010011111100",
								"0001001111100010",
								"0001000100001110",
								"1110000000001010",
								"1001010100001110",
								"1011111101010010",
								"1101110100001111",
								"1101000111011101",
								"1111000011000110",
								"1110001100101001",
								"1111011110111111",
								"1110110011110111",
								"1111101000010100",
								"1111001011000010",
								"1111101100010001",
								"1111011000110010",
								"1111101100000111",
								"1111011101000110",
								"1111101010001010",
								"1111100011100101",
								"1111101010111011",
								"1111100111111001",
								"1111101010111100",
								"1111101010110100",
								"1111101100010001",
								"1111101101000101",
								"1111101011101111",
								"1111101110111111",
								"1111101101100010",
								"1111110000000010",
								"1111101110000101",
								"1111110001001011",
								"1111101111000100",
								"1111110010010001",
								"1111101111110001",
								"1111110011011110",
								"1111110000100110",
								"1111110011111101",
								"1111110001110001",
								"1111110100001010",
								"1111110010000110",
								"1111110101010001",
								"1111110010111111",
								"1111110100111110",
								"1111110110011110",
								"0001011000010001",
								"0101101001001001",
								"0101111001000011",
								"0011011110011101",
								"0100011010100000",
								"0010111111000100",
								"0011010101001011",
								"0010101011111010",
								"0010101111011101",
								"0010011101000100",
								"0010010100110011",
								"0010010000010000",
								"0010000011101000",
								"0010000101101010",
								"0001111000001100",
								"0001111100100110",
								"0001101100010100",
								"0001110010111000",
								"0001100101110110",
								"0001101101100011",
								"0001100001111000",
								"0001101001011011",
								"0001011110000100",
								"0001100101111010",
								"0001011011011111",
								"0001100010000000",
								"0001011000110101",
								"0001011111101010",
								"0001010110010011",
								"0001011101001100",
								"0001010100001100",
								"0001011010110000",
								"0001010010100110",
								"0001011000100111",
								"0001010001000011",
								"0001010110011110",
								"0001001111100000",
								"0001010100010100",
								"0001001110000100",
								"0001010010110101",
								"0001001101010110",
								"0000110000000010",
								"1100101100110011",
								"1001001001110111",
								"1100111011010010",
								"1101010111111101",
								"1101100100111110",
								"1110110111001110",
								"1110001111001110",
								"1111011010010010",
								"1110101100010000",
								"1111101001011011",
								"1111000100001110",
								"1111110001110111",
								"1111001111111011",
								"1111110100001110",
								"1111011000100100",
								"1111110011110100",
								"1111011110100010",
								"1111110011000110",
								"1111011111001111",
								"1111101111101001",
								"1111100010100110",
								"1111110000100111",
								"1111100100111110",
								"1111101111111001",
								"1111100111011011",
								"1111110000111101",
								"1111101001000000",
								"1111110000100110",
								"1111101010000110",
								"1111110010001000",
								"1111101011011000",
								"1111110001111100",
								"1111101100101100",
								"1111110010100010",
								"1111101101110011",
								"1111110010100111",
								"1111101110111100",
								"1111110011000101",
								"1111101111100011",
								"1111110011110111",
								"1111101111110001",
								"1111111101101011",
								"0010001001101010",
								"0110010111111011",
								"0101000110001101",
								"0011100111000110",
								"0100001111000101",
								"0010110101011001",
								"0011010110010010",
								"0010011100110111",
								"0010101111001011",
								"0010001100011001",
								"0010010100110000",
								"0010000010011110",
								"0010000111011110",
								"0001111100111011",
								"0001111010110110",
								"0001110110101000",
								"0001110010001000",
								"0001110001000111",
								"0001101011000100",
								"0001101011111111",
								"0001100010110100",
								"0001100100100011",
								"0001011101101101",
								"0001100001010000",
								"0001011010101010",
								"0001011110101110",
								"0001011000010010",
								"0001011100001001",
								"0001010101110000",
								"0001011001001001",
								"0001010011001010",
								"0001010111100100",
								"0001010001110010",
								"0001010101000011",
								"0001001111100111",
								"0001010011100100",
								"0001001110000111",
								"0001010001001011",
								"0001001100111011",
								"0001001111111000",
								"0001001010111111",
								"0000001110011101",
								"1011011000010001",
								"1001011111011110",
								"1101100111011110",
								"1100111100110000",
								"1110001000110101",
								"1110100001100010",
								"1110100010110011",
								"1111001101100101",
								"1110110101000111",
								"1111100000100001",
								"1111000010000111",
								"1111101001100100",
								"1111001010100111",
								"1111101110011010",
								"1111010101110011",
								"1111110100011011",
								"1111011010001011",
								"1111110101001110",
								"1111011110001001",
								"1111110101011001",
								"1111100001010000",
								"1111110100101101",
								"1111100001001011",
								"1111110000110110",
								"1111100010010100",
								"1111110001101010",
								"1111100011101101",
								"1111110001101001",
								"1111100101111001",
								"1111110010010011",
								"1111100111000000",
								"1111110010000110",
								"1111100111010010",
								"1111110011100100",
								"1111101001000001",
								"1111110011001110",
								"1111101001100001",
								"1111110011001010",
								"1111101011100011",
								"1111110010111110",
								"1111101011110011",
								"0000001001110111",
								"0011000101000001",
								"0110101110001000",
								"0100010011101111",
								"0011111001010011",
								"0011110111110101",
								"0010110110110001",
								"0011001110100001",
								"0010010110110001",
								"0010101101100010",
								"0010000100011111",
								"0010010101101111",
								"0001111000010111",
								"0010000100101110",
								"0001110000011011",
								"0001111000101100",
								"0001101011011100",
								"0001110011011111",
								"0001101010110001",
								"0001101100101110",
								"0001100110111000",
								"0001100111111001",
								"0001100011011100",
								"0001100011010101",
								"0001011111111000",
								"0001011101000110",
								"0001011000101001",
								"0001011000100110",
								"0001010111001011",
								"0001010110001111",
								"0001010100001101",
								"0001010011111111",
								"0001010010101010",
								"0001010001111101",
								"0001010000101001",
								"0001001111000001",
								"0001001111011111",
								"0001001101101110",
								"0001001100111110",
								"0001001100010101",
								"0001001100000100",
								"0001001000000001",
								"1111011100000110",
								"1010001101011011",
								"1010010000111001");
								
	variable expected_out : WAV_IN := ("0000000000011101",
										"1111111111010001",
										"1111111011010011",
										"1111110110111010",
										"1111110010110000",
										"1111101111000011",
										"1111101111010010",
										"1111101111110111",
										"1111101111100010",
										"1111110001010101",
										"1111110100111100",
										"1111111001011011",
										"1111111101100011",
										"0000000001011100",
										"1111111111010000",
										"1111111011100011",
										"1111110101010001",
										"1111101100100010",
										"1111100101110110",
										"1111011111100110",
										"1111011010110100",
										"1111010101010111",
										"1111010001100001",
										"1111001100010011",
										"1111001000011101",
										"1111000101111001",
										"1111000010010001",
										"1110111111010001",
										"1110111011110100",
										"1110111000101000",
										"1110110101110100",
										"1110110010111001",
										"1110110000010110",
										"1110101101110111",
										"1110101100010111",
										"1110101011010000",
										"1110101000000110",
										"1110100110000011",
										"1110100010101010",
										"1110011111000000",
										"1110011101010001",
										"1110011010101110",
										"1110011000100111",
										"1110010110001101",
										"1110010100001101",
										"1110010000111101",
										"1110001010011000",
										"1110000011010110",
										"1101111101011100",
										"1101110111011111",
										"1101110101000010",
										"1101110011100111",
										"1101110001100001",
										"1101110000110101",
										"1101110001111111",
										"1101110101000011",
										"1101110110111101",
										"1101111000110100",
										"1101110111100011",
										"1101110100111010",
										"1101110011010110",
										"1101110001011111",
										"1101110000101010",
										"1101110000001000",
										"1101101111001011",
										"1101101101010100",
										"1101101100000101",
										"1101101010010000",
										"1101101000010000",
										"1101100111000011",
										"1101100101101001",
										"1101100011101010",
										"1101100010001011",
										"1101100000101010",
										"1101011110111110",
										"1101011110000100",
										"1101011111001001",
										"1101100100011001",
										"1101100111110111",
										"1101101011000110",
										"1101101100011000",
										"1101101001101011",
										"1101101000110101",
										"1101100111110010",
										"1101100111001110",
										"1101100111000010",
										"1101100110111110",
										"1101100111010010",
										"1101100110111011",
										"1101100101101010",
										"1101100001011111",
										"1101011100110100",
										"1101011001000100",
										"1101010101110011",
										"1101010110001101",
										"1101010111000001",
										"1101010111011111",
										"1101011001001100",
										"1101011100001100",
										"1101100001000100",
										"1101100110100000",
										"1101101010110111",
										"1101101101000100",
										"1101101110110001",
										"1101101110001111",
										"1101101111101000",
										"1101110000001110",
										"1101110001101001",
										"1101110011010011",
										"1101110011100001",
										"1101110101001000",
										"1101110100101011",
										"1101110101100101",
										"1101110110100110",
										"1101110111001101",
										"1101110111111111",
										"1101111000011100",
										"1101110111111000",
										"1101100010111111",
										"1100101001110111",
										"1011111010111011",
										"1011011000011000",
										"1011000011100000",
										"1011011110101111",
										"1011101001101100",
										"1011110001000011",
										"1011111011010010",
										"1011111110010010",
										"1100000101001011",
										"1100000111000110",
										"1100001011000001",
										"1100001100001000",
										"1100001110010100",
										"1100001110000111",
										"1100001011101100",
										"1100000110100111",
										"1100000011001101",
										"1011111110111000",
										"1011111110001000",
										"1011111110011010",
										"1011111110100010",
										"1011111111000000",
										"1100000001101101",
										"1100000110000111",
										"1100001010000111",
										"1100001110010101",
										"1100001111101011",
										"1100001110110100",
										"1100001110010011",
										"1100001101001100",
										"1100001100110010",
										"1100001101001110",
										"1100001101010101",
										"1100001100011101",
										"1100001100101110",
										"1100001011111001",
										"1100001011000100",
										"1100001010111000",
										"1100001010111001",
										"1100100011000100",
										"1110101100000101",
										"0001100010010000",
										"0010111001101111",
										"0100001010100001",
										"0011001110000000",
										"0001011101101110",
										"0001001001010001",
										"0000010110010001",
										"0000000110110101",
										"1111110000111101",
										"1111100110100010",
										"1111011101000010",
										"1111010101111011",
										"1111010001010101",
										"1111001100101100",
										"1111001010110011",
										"1111000111011110",
										"1111000110010110",
										"1111000000000101",
										"1110111010101010",
										"1110110100111000",
										"1110110000111100",
										"1110101101110111",
										"1110101111000110",
										"1110101101010110",
										"1110101110101101",
										"1110110000010000",
										"1110110100111110",
										"1110110111111111",
										"1110111100000001",
										"1110111101110011",
										"1110111101101100",
										"1110111101101001",
										"1110111100111100",
										"1110111100001101",
										"1110111101001101",
										"1110111101010101",
										"1110111101110000",
										"1110111110000000",
										"1110111101100101",
										"1110111101001001",
										"1110110001110101",
										"1101000111100001",
										"1001111110001110",
										"0111111011001101",
										"0110001011011010",
										"0101111011111001",
										"0111100111011000",
										"1000000000011011",
										"1000101100010011",
										"1001001000111000",
										"1001011110010011",
										"1001110100011011",
										"1010000000111100",
										"1010010000011011",
										"1010010111110000",
										"1010100011000111",
										"1010100111010101",
										"1010101111101011",
										"1010110011000010",
										"1010111000101011",
										"1010111010111100",
										"1010111011100011",
										"1010110111110000",
										"1010110110011001",
										"1010110011101101",
										"1010110100001110",
										"1010110111001100",
										"1010111000100000",
										"1010111001111101",
										"1010111101111111",
										"1011000011000011",
										"1011001000100101",
										"1011001101011000",
										"1011010000111001",
										"1011010001100110",
										"1011010010101110",
										"1011010011010101",
										"1011010011110000",
										"1011010100111001",
										"1011010110101101",
										"1011010110101111",
										"1011011010100000",
										"1100110001010010",
										"0010000011100001",
										"0111010010100111",
										"1001110010001001",
										"1011110010110001",
										"1000011110111001",
										"0101100011001111",
										"0100110001001011",
										"0011001001001110",
										"0010110010000111",
										"0001111101011110",
										"0001101111101110",
										"0001010101010101",
										"0001001011111111",
										"0000111110011001",
										"0000110111101100",
										"0000101111111001",
										"0000101011011110",
										"0000100110101010",
										"0000100010110110",
										"0000011111111100",
										"0000011100001101",
										"0000011010100001",
										"0000010100100000",
										"0000001101100100",
										"0000000110010101",
										"0000000000011111",
										"1111111100000010",
										"1111111100001010",
										"1111111001110001",
										"1111111001101010",
										"1111111001111001",
										"1111111101011101",
										"0000000000110100",
										"0000000011110111",
										"0000000100101010",
										"0000000100000001",
										"0000000001111111",
										"0000000001111100",
										"0000000000100111",
										"0000000000100001",
										"0000000000000111",
										"1111011100000000",
										"1100001001010111",
										"0111010001010110",
										"0100010111101001",
										"0001101101111100",
										"0010010011100000",
										"0100110010101101",
										"0101010001011010",
										"0110100001110011",
										"0111000100000011",
										"0111101110111110",
										"1000001011100111",
										"1000100011101000",
										"1000111001010111",
										"1001000111111110",
										"1001010111101000",
										"1001100001011010",
										"1001101101100110",
										"1001110100010111",
										"1001111101010000",
										"1010000010010011",
										"1010001000110110",
										"1010001100100101",
										"1010010010000010",
										"1010010100001100",
										"1010010110001110",
										"1010010011001110",
										"1010010010001011",
										"1010010000010100",
										"1010010000110011",
										"1010010011101100",
										"1010010110001100",
										"1010011000100001",
										"1010011100110100",
										"1010100010100010",
										"1010101001100111",
										"1010101110101110",
										"1010110011100000",
										"1010110100010110",
										"1010110110001100",
										"1010110110111010",
										"1011000000111111",
										"1101100110101000",
										"0100111100110000",
										"1010011110011000",
										"1101100010010011",
										"1111000001001011",
										"1001111001100110",
										"0111010110000100",
										"0110000010100101",
										"0100010100111111",
										"0011110111011000",
										"0010111000100111",
										"0010101100000011",
										"0010000111101100",
										"0010000001100001",
										"0001101100011001",
										"0001101000101101",
										"0001011100000111",
										"0001011001001000",
										"0001010000101001",
										"0001001110011010",
										"0001001000000111",
										"0001000110001010",
										"0001000001101010",
										"0000111111011100",
										"0000111100011111",
										"0000111001100011",
										"0000110111010010",
										"0000110011000001",
										"0000101011100011",
										"0000100100111111",
										"0000011110101110",
										"0000011001110010",
										"0000011000110110",
										"0000010111101010",
										"0000010110001010",
										"0000010110000101",
										"0000011001000100",
										"0000011011001100",
										"0000011110101110",
										"0000100000010101",
										"0000100000010000",
										"0000011101100100",
										"1111010000100000",
										"1010001101000101",
										"0100011111101011",
										"0001001010110101",
										"1110001101000000",
										"0000010000000001",
										"0010110100011010",
										"0011011110101101",
										"0101000110110011",
										"0101101010100001",
										"0110100111101011",
										"0111000100001110",
										"0111101010010010",
										"1000000000001101",
										"1000011000101011",
										"1000101001111000",
										"1000111001100011",
										"1001000111001100",
										"1001010010001111",
										"1001011100110110",
										"1001100101010100",
										"1001101101110100",
										"1001110100010010",
										"1001111011010111",
										"1010000000100111",
										"1010000110100101",
										"1010001010111000",
										"1010010000010100",
										"1010010011101010",
										"1010010110101011",
										"1010010101011111",
										"1010010100101011",
										"1010010011011010",
										"1010010011100110",
										"1010010111000100",
										"1010011010000011",
										"1010011100111001",
										"1010100001010110",
										"1010100111011000",
										"1010101111011110",
										"1010110101010001",
										"1011010100000000",
										"1111001110111101",
										"0111001100010100",
										"1011101101110111",
										"1110111110100111",
										"1110110011001101",
										"1001001001111000",
										"0111100110010001",
										"0101110000000010",
										"0100011110110110",
										"0011110011010111",
										"0010111101101110",
										"0010101110011000",
										"0010001100101110",
										"0010000110000100",
										"0001110001000101",
										"0001101110010011",
										"0001011111000000",
										"0001011110010001",
										"0001010100000011",
										"0001010010111000",
										"0001001011011011",
										"0001001010011111",
										"0001000011110101",
										"0001000011000110",
										"0000111110000110",
										"0000111101001000",
										"0000111001011011",
										"0000111000010011",
										"0000110100110000",
										"0000110011110101",
										"0000110000101001",
										"0000101101110000",
										"0000100110110011",
										"0000100000001100",
										"0000011010010111",
										"0000010101001111",
										"0000010011101111",
										"0000010010110000",
										"0000010000110000",
										"0000010001010000",
										"0000010011000001",
										"0000010000100000",
										"1110010101001101",
										"1000011001000100",
										"0011001000100100",
										"1111101101100000",
										"1101011010001100",
										"0000100000101010",
										"0010011001011001",
										"0011011000000010",
										"0100111000011000",
										"0101011100001101",
										"0110011100001001",
										"0110110101011101",
										"0111011110010100",
										"0111110001110110",
										"1000001101010011",
										"1000011100000101",
										"1000101111010111",
										"1000111011001000",
										"1001001000011001",
										"1001010001011010",
										"1001011011010101",
										"1001100011000100",
										"1001101010101111",
										"1001110001001001",
										"1001110111011101",
										"1001111100101011",
										"1010000010001001",
										"1010000111001001",
										"1010001011100100",
										"1010001111111010",
										"1010010011100000",
										"1010010111110111",
										"1010011011000000",
										"1010011101011000",
										"1010011100010011",
										"1010011010011111",
										"1010011001000010",
										"1010011001001100",
										"1010011011010011",
										"1010011110110100",
										"1010100001001000",
										"1011010110110000",
										"0000101011000010",
										"1000100100011001",
										"1100010101110110",
										"1111101101001101",
										"1101101010100001",
										"1000011001000000",
										"0111011001100110",
										"0101001101110000",
										"0100011001001111",
										"0011011111111011",
										"0010111011110010",
										"0010100011001011",
										"0010001010011111",
										"0010000000000000",
										"0001101101110010",
										"0001101001101111",
										"0001011101001000",
										"0001011011001110",
										"0001010001100010",
										"0001010000101101",
										"0001001000110001",
										"0001000111110010",
										"0001000010001110",
										"0001000001010100",
										"0000111101000000",
										"0000111100001110",
										"0000110111011100",
										"0000110111000110",
										"0000110011001101",
										"0000110010011001",
										"0000101111110000",
										"0000101110011000",
										"0000101011010011",
										"0000101011000010",
										"0000101000011010",
										"0000100110111111",
										"0000100000101000",
										"0000011010101000",
										"0000010011110111",
										"0000001111001110",
										"0000001101001110",
										"1111111100110110",
										"1101000000011011",
										"0110011100111111",
										"0001110101001110",
										"1110010100011111",
										"1101001011010111",
										"0000111001100000",
										"0010001000111111",
										"0011100000010001",
										"0100101110110010",
										"0101011010011011",
										"0110010100010000",
										"0110110000000111",
										"0111011000110110",
										"0111101011011001",
										"1000001000001100",
										"1000010100111110",
										"1000101001000101",
										"1000110011101010",
										"1001000010011001",
										"1001001010111111",
										"1001010110001000",
										"1001011101000111",
										"1001100101101111",
										"1001101011011101",
										"1001110010101110",
										"1001110111111110",
										"1001111101111111",
										"1010000010001111",
										"1010000111010000",
										"1010001011010101",
										"1010001111011000",
										"1010010011100001",
										"1010010111011110",
										"1010011010110010",
										"1010011110110000",
										"1010100001111101",
										"1010100100111011",
										"1010100111011010",
										"1010100110000111",
										"1010100011100000",
										"1010100100101100",
										"1011111111111000",
										"0010100010010000",
										"1001101100000001",
										"1100111011000000",
										"1111110110010100",
										"1100000001101101",
										"0111110110010011",
										"0110111111000010",
										"0100110100101111",
										"0100010101001111",
										"0011010000001010",
										"0010111010110111",
										"0010011001000100",
										"0010001010001101",
										"0001111001101001",
										"0001101111110000",
										"0001100110111011",
										"0001011111001110",
										"0001011001111110",
										"0001010010101011",
										"0001010000000110",
										"0001001010010100",
										"0001001000011011",
										"0001000011000000",
										"0001000001101100",
										"0000111101011101",
										"0000111100011111",
										"0000111000110010",
										"0000111000000101",
										"0000110100100100",
										"0000110011100111",
										"0000110000111011",
										"0000101111011100",
										"0000101101000101",
										"0000101100011101",
										"0000101001100110",
										"0000101001011000",
										"0000100110110111",
										"0000100110001000",
										"0000100100001110",
										"0000100010111100",
										"0000011110000000",
										"1111110011111101",
										"1011101011111000",
										"0100111001000111",
										"0000110010100111",
										"1101001010000100",
										"1101011010110101",
										"0001000100001100",
										"0001111000100011",
										"0011101001011110",
										"0100100110101011",
										"0101100100000011",
										"0110010100001110",
										"0110110100111010",
										"0111011000000101",
										"0111101100111001",
										"1000000110001101",
										"1000010101001111",
										"1000101001001111",
										"1000110011101001",
										"1001000011010100",
										"1001001011011111",
										"1001010110000101",
										"1001011101011000",
										"1001100110000001",
										"1001101011111100",
										"1001110011011101",
										"1001111000000110",
										"1001111110110111",
										"1010000010110101",
										"1010001000110100",
										"1010001100011011",
										"1010010001100000",
										"1010010101000011",
										"1010011001011100",
										"1010011100110001",
										"1010100000100011",
										"1010100011101111",
										"1010100111011100",
										"1010101011000000",
										"1010101110001101",
										"1010110000011001",
										"1010111001011111",
										"1101001111100000",
										"0100101100001011",
										"1010110011000101",
										"1101111000110011",
										"1111110110010010",
										"1010101100110001",
										"0111100111101110",
										"0110011001010111",
										"0100011011010010",
										"0100000001010100",
										"0011000000010011",
										"0010110111011011",
										"0010010101010101",
										"0010001110111111",
										"0001111001000011",
										"0001110100000010",
										"0001100110110110",
										"0001100010110111",
										"0001011010111001",
										"0001011000000100",
										"0001010010000001",
										"0001001111000001",
										"0001001011111100",
										"0001000111001111",
										"0001000110000001",
										"0001000011010000",
										"0001000000011010",
										"0000111110100100",
										"0000111100011100",
										"0000111001101011",
										"0000111000100011",
										"0000110110011010",
										"0000110100100111",
										"0000110010111100",
										"0000110001011100",
										"0000101110111101",
										"0000101110100011",
										"0000101100010011",
										"0000101011100011",
										"0000101001110111",
										"0000101001001010",
										"0000100110110110",
										"1111101001000101",
										"1010101010011110",
										"0100001000011010",
										"0000010100010101",
										"1100101110110000",
										"1110001011000110",
										"0001010100111111",
										"0001111111100001",
										"0011110011101100",
										"0100011111010110",
										"0101100001010011",
										"0110000111111100",
										"0110110011011011",
										"0111010100111011",
										"0111110001110111",
										"1000001011101000",
										"1000011100000011",
										"1000101101110111",
										"1000111000110000",
										"1001000101101100",
										"1001001110110111",
										"1001011010100010",
										"1001100010000100",
										"1001101011000000",
										"1001110001010010",
										"1001110111010110",
										"1001111100111110",
										"1010000011011111",
										"1010000111100011",
										"1010001101101001",
										"1010010001100010",
										"1010010110101000",
										"1010011001111111",
										"1010011110111011",
										"1010100001110110",
										"1010100110010111",
										"1010101001111110",
										"1010101101011101",
										"1010110000010001",
										"1010110011111010",
										"1010110101111111",
										"1011000111101011",
										"1110011000001010",
										"0110010111111000",
										"1011101010001000",
										"1110111010000111",
										"1111110010110100",
										"1010000011111100",
										"0111110100100101",
										"0110001001110101",
										"0100011101011011",
										"0011111000001101",
										"0010111001110100",
										"0010101100100010",
										"0010000111100111",
										"0010000011110100",
										"0001110001110000",
										"0001110011110111",
										"0001101001000100",
										"0001101010010000",
										"0001011111011101",
										"0001011110101011",
										"0001010111011100",
										"0001010110000110",
										"0001010000111010",
										"0001010000000111",
										"0001001011111100",
										"0001001010101011",
										"0001000111101110",
										"0001000101011000",
										"0001000011001100",
										"0001000001101010",
										"0000111111011011",
										"0000111101101111",
										"0000111011011100",
										"0000111001111010",
										"0000111000001110",
										"0000110110001110",
										"0000110101100010",
										"0000110100000010",
										"0000110010101110",
										"0000110001100000",
										"0000110000101100",
										"0000101100010100",
										"1111001001010100",
										"1001010011001010",
										"0011001111000101",
										"1111100111000110",
										"1100100100110111",
										"1111001110111100",
										"0001110010110100",
										"0010100101010111",
										"0100010000011010",
										"0100110010011010",
										"0101110010110010",
										"0110001110011100",
										"0110111010010001",
										"0111010001101011",
										"0111101110010010",
										"1000000001111100",
										"1000011001010000",
										"1000101100000010",
										"1000111110011000",
										"1001001101011011",
										"1001010111110111",
										"1001100001010100",
										"1001101001000110",
										"1001110000101111",
										"1001110111001000",
										"1001111110100011",
										"1010000011110010",
										"1010001010000010",
										"1010001111001110",
										"1010010100000010",
										"1010011000101011",
										"1010011101100101",
										"1010100001010010",
										"1010100101110111",
										"1010101001000000",
										"1010101101010010",
										"1010110000011000",
										"1010110100101011",
										"1010110111101010",
										"1010111011010011",
										"1010111101011101",
										"1011100001101111",
										"0000000011000000",
										"1000001011111110",
										"1100011110000010",
										"1111110110000111",
										"1110111101111100",
										"1001010000100101",
										"0111111100101001",
										"0101111010010100",
										"0100110011000010",
										"0100000000110101",
										"0011001011110101",
										"0010110100010000",
										"0010010000100101",
										"0010000101110010",
										"0001110001011100",
										"0001101111011111",
										"0001100000111000",
										"0001100010000000",
										"0001011011010101",
										"0001011111100000",
										"0001011011011100",
										"0001011101111011",
										"0001011000001100",
										"0001010111111100",
										"0001010011000111",
										"0001010010110001",
										"0001001110101111",
										"0001001110000010",
										"0001001011010111",
										"0001001010001100",
										"0001000111110100",
										"0001000110011110",
										"0001000011111000",
										"0001000011011110",
										"0001000001000011",
										"0001000000011000",
										"0000111110001000",
										"0000111101100101",
										"0000111011110101",
										"0000111010100101",
										"0000111001110000",
										"0000101111001010",
										"1110010101000011",
										"0111110000111111",
										"0010011010100011",
										"1110110001001000",
										"1100101011101101",
										"0000001110001111",
										"0001111110001010",
										"0011001000011001",
										"0100101000010011",
										"0101010001010011",
										"0110010010110101",
										"0110101101001110",
										"0111010100111011",
										"0111100100011001",
										"0111111110010011",
										"1000001010001001",
										"1000011111011111",
										"1000101011010011",
										"1000111011000101",
										"1001000101101110",
										"1001010101000010",
										"1001100001100110",
										"1001101110111101",
										"1001111001101100",
										"1010000001110110",
										"1010000111101011",
										"1010001101000110",
										"1010010010001101",
										"1010010111000111",
										"1010011100101100",
										"1010100001110100",
										"1010100110011001",
										"1010101010010111",
										"1010101110011101",
										"1010110010000000",
										"1010110110000000",
										"1010111001101011",
										"1010111101100011",
										"1011000000001111",
										"1011000011111011",
										"1011000111000011",
										"1100001001110001",
										"0001111110011011",
										"1001101110110101",
										"1101010010010110",
										"0000100100000011",
										"1101110011011111",
										"1000110001011011",
										"0111110110000110",
										"0101100101010001",
										"0100111000111111",
										"0011111010000000",
										"0011011010101100",
										"0010111110101101",
										"0010101001001101",
										"0010011011010100",
										"0010000111101000",
										"0001111100110001",
										"0001101101001101",
										"0001100110011001",
										"0001011110000011",
										"0001011101000101",
										"0001010110000000",
										"0001010110100001",
										"0001010011011111",
										"0001011000000010",
										"0001010110111110",
										"0001011010000001",
										"0001010111011111",
										"0001010110101100",
										"0001010011000111",
										"0001010010011110",
										"0001001111001011",
										"0001001110101110",
										"0001001101010101",
										"0001001100000100",
										"0001001010000011",
										"0001001000111011",
										"0001000110101100",
										"0001000111000110",
										"0001000100100100",
										"0001000100110100",
										"0001000010100010",
										"0000101011110101",
										"1101010010010111",
										"0110010111001101",
										"0001101111010001",
										"1101111111110101",
										"1101001101000001",
										"0001000100011000",
										"0010001001100110",
										"0011101100001000",
										"0100110110011011",
										"0101101000101101",
										"0110100001011111",
										"0110111111111001",
										"0111101000101101",
										"0111111100110001",
										"1000011001110100",
										"1000100110101111",
										"1000110111111110",
										"1000111101101000",
										"1001001001100110",
										"1001001110001010",
										"1001011001110000",
										"1001100001000101",
										"1001101010011110",
										"1001110001011110",
										"1001111100010001",
										"1010000111000100",
										"1010010001110011",
										"1010011010100000",
										"1010100001010111",
										"1010100101110011",
										"1010101010011010",
										"1010101110111011",
										"1010110011001101",
										"1010110110110001",
										"1010111011101111",
										"1010111110111010",
										"1011000011001001",
										"1011000110110100",
										"1011001001100000",
										"1011001100111011",
										"1011010010101000",
										"1101000011100000",
										"0100000010011010",
										"1010111101100101");
	
	
	begin
		
		-- inital reset of the filter
		rst_l <= '0';
		wait until clk'event and clk='1';
		rst_l <= '1'; 
		
		-- loop over all the samples
		for i in 0 to SAMPLES-1 loop	
			
			sample <= input(i);
			expected <= expected_out(i);
			
			
			wait until clk'event and clk='1'; 
			
			-- If the actual output and the expected output
			-- mismatch, raise an asserion
			assert (output = expected)
			report "Mismatch for index i = " & integer'image(i)
			severity error;
			
		end loop;	 
		
		enable <= '0';
		end process;

end TB_Arch;

