library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all; 

entity IIR_TB_Street is
end IIR_TB_Street;

architecture TB_Arch of IIR_TB_Street is	

component IIR  
	generic (Nbit : natural := 8);
	port (
		clk		:	in	std_logic;
		rst_l	:	in	std_logic;
		x		:	in	std_logic_vector(Nbit-1 downto 0);	
		y		:	out	std_logic_vector(Nbit-1 downto 0)
	);
end component;

	constant BITS		:	natural	:=	16;
	constant SAMPLES 	:	natural	:= 	1000;

	signal clk		: 	std_logic	:= '0'; 
	signal rst_l 	: 	std_logic;
	signal sample	:	std_logic_vector(BITS-1 downto 0);
	signal output	:	std_logic_vector(BITS-1 downto 0);
	signal expected	:	std_logic_vector(BITS-1 downto 0);
	
	signal enable	:	std_logic	:=	'1';
	
	type WAV_IN is array (0 to SAMPLES-1) of std_logic_vector(BITS-1 downto 0);

begin
	
	filter: IIR
	generic map(BITS)
	port map(clk, rst_l, sample, output);
	
	clk <= not clk and enable after 11338 ns; -- 44100Hz clock
	
	driver_p: process
	
	variable input : WAV_IN := ("1111111100110100",
								"1111111100011000",
								"1111111101000000",
								"1111111100111001",
								"1111111101001100",
								"1111111100110010",
								"1111111100101011",
								"1111111100000001",
								"1111111011101110",
								"1111111011001001",
								"1111111011001110",
								"1111111011001000",
								"1111111011101000",
								"1111111100001011",
								"1111111100111110",
								"1111111101100110",
								"1111111110010010",
								"1111111110101100",
								"1111111111000000",
								"1111111111000001",
								"1111111111000111",
								"1111111111000010",
								"1111111111000111",
								"1111111111001000",
								"1111111111011101",
								"1111111111111000",
								"0000000000011011",
								"0000000000111111",
								"0000000001101000",
								"0000000010001011",
								"0000000010100010",
								"0000000010110110",
								"0000000010111110",
								"0000000010111110",
								"0000000010111001",
								"0000000010100110",
								"0000000010010011",
								"0000000001111100",
								"0000000001100111",
								"0000000001100111",
								"0000000001100000",
								"0000000001110001",
								"0000000001101111",
								"0000000001111100",
								"0000000001111000",
								"0000000001110000",
								"0000000001100010",
								"0000000001010000",
								"0000000001000000",
								"0000000000111001",
								"0000000000111101",
								"0000000001001010",
								"0000000001100010",
								"0000000010000110",
								"0000000010011110",
								"0000000010110101",
								"0000000010111001",
								"0000000010110011",
								"0000000010101010",
								"0000000010000100",
								"0000000001100100",
								"0000000000110001",
								"0000000000001100",
								"1111111111011101",
								"1111111111000000",
								"1111111110110001",
								"1111111110110010",
								"1111111111000001",
								"1111111111011010",
								"1111111111110101",
								"0000000000001111",
								"0000000000110001",
								"0000000000111101",
								"0000000001000110",
								"0000000000110111",
								"0000000000011101",
								"1111111111111111",
								"1111111111011001",
								"1111111110111101",
								"1111111110101010",
								"1111111110011010",
								"1111111110011010",
								"1111111110010101",
								"1111111110010101",
								"1111111110010101",
								"1111111110010100",
								"1111111110011101",
								"1111111110100101",
								"1111111110110110",
								"1111111111000010",
								"1111111111011010",
								"1111111111100101",
								"1111111111101110",
								"1111111111110000",
								"1111111111101001",
								"1111111111100010",
								"1111111111010100",
								"1111111111010000",
								"1111111111001111",
								"1111111111001110",
								"1111111111011011",
								"1111111111100100",
								"1111111111111000",
								"1111111111111011",
								"1111111111111011",
								"1111111111101110",
								"1111111111011100",
								"1111111111000101",
								"1111111110101011",
								"1111111110011110",
								"1111111110001100",
								"1111111110001010",
								"1111111110000011",
								"1111111110000100",
								"1111111110000010",
								"1111111110010001",
								"1111111110011101",
								"1111111110110001",
								"1111111110111111",
								"1111111111001011",
								"1111111111010111",
								"1111111111010010",
								"1111111111010010",
								"1111111110111110",
								"1111111110110011",
								"1111111110011101",
								"1111111110011010",
								"1111111110010011",
								"1111111110011000",
								"1111111110010111",
								"1111111110100101",
								"1111111110011011",
								"1111111110011111",
								"1111111110100011",
								"1111111110101101",
								"1111111110111100",
								"1111111111000101",
								"1111111111010000",
								"1111111111000100",
								"1111111110111101",
								"1111111110100010",
								"1111111110010101",
								"1111111110000010",
								"1111111110000000",
								"1111111110000100",
								"1111111110010110",
								"1111111110101010",
								"1111111110111001",
								"1111111111001000",
								"1111111111001011",
								"1111111111010010",
								"1111111111011011",
								"1111111111100110",
								"1111111111111101",
								"0000000000011101",
								"0000000000111110",
								"0000000001011011",
								"0000000001111000",
								"0000000010000111",
								"0000000010011001",
								"0000000010101000",
								"0000000010011111",
								"0000000010010110",
								"0000000010000001",
								"0000000010000000",
								"0000000001110111",
								"0000000010001100",
								"0000000010011010",
								"0000000010110100",
								"0000000011000111",
								"0000000011011000",
								"0000000011011001",
								"0000000011010101",
								"0000000011000011",
								"0000000010100001",
								"0000000001110010",
								"0000000000110111",
								"0000000000000010",
								"1111111111010111",
								"1111111110111100",
								"1111111110101110",
								"1111111111000011",
								"1111111111010100",
								"1111111111111001",
								"0000000000011000",
								"0000000000110010",
								"0000000001000100",
								"0000000001001100",
								"0000000001001110",
								"0000000001010000",
								"0000000001011001",
								"0000000001011001",
								"0000000001010010",
								"0000000001001001",
								"0000000000101110",
								"0000000000010010",
								"1111111111110111",
								"1111111111011110",
								"1111111110111110",
								"1111111110100101",
								"1111111110011010",
								"1111111110100100",
								"1111111111000010",
								"1111111111101000",
								"0000000000000011",
								"0000000000000101",
								"1111111111111111",
								"1111111111101110",
								"1111111111011000",
								"1111111110110000",
								"1111111110000010",
								"1111111101001100",
								"1111111100001110",
								"1111111011011101",
								"1111111010101010",
								"1111111010011111",
								"1111111010110111",
								"1111111011100011",
								"1111111100110001",
								"1111111101100011",
								"1111111110100010",
								"1111111110101011",
								"1111111110110011",
								"1111111110011010",
								"1111111110000010",
								"1111111101110110",
								"1111111101111110",
								"1111111110100101",
								"1111111111100000",
								"0000000000000101",
								"0000000000101001",
								"0000000000101011",
								"0000000000011110",
								"0000000000100001",
								"0000000000001011",
								"0000000000001011",
								"0000000000000001",
								"0000000000000101",
								"0000000000010010",
								"0000000000001111",
								"0000000000100101",
								"0000000000101101",
								"0000000000111001",
								"0000000000111010",
								"0000000000110111",
								"0000000000110110",
								"0000000000110000",
								"0000000000101010",
								"0000000000100100",
								"0000000000100010",
								"0000000000011000",
								"0000000000001110",
								"0000000000000110",
								"1111111111111100",
								"1111111111101111",
								"1111111111010111",
								"1111111111001100",
								"1111111110110111",
								"1111111110111100",
								"1111111110111011",
								"1111111111011010",
								"1111111111101110",
								"0000000000001111",
								"0000000000010011",
								"0000000000001110",
								"1111111111111101",
								"1111111111011100",
								"1111111110111011",
								"1111111110101100",
								"1111111110011101",
								"1111111110101011",
								"1111111110111111",
								"1111111111011101",
								"1111111111110101",
								"0000000000000010",
								"1111111111111110",
								"1111111111110010",
								"1111111111010100",
								"1111111110101001",
								"1111111101111001",
								"1111111101000011",
								"1111111100010101",
								"1111111100000010",
								"1111111011111100",
								"1111111100011110",
								"1111111101001100",
								"1111111110010001",
								"1111111111010101",
								"0000000000001100",
								"0000000000110001",
								"0000000001001111",
								"0000000001010101",
								"0000000001011011",
								"0000000001100100",
								"0000000001110010",
								"0000000010001001",
								"0000000010100010",
								"0000000011000011",
								"0000000011100101",
								"0000000011111000",
								"0000000100011000",
								"0000000100100111",
								"0000000100110000",
								"0000000100101010",
								"0000000100011100",
								"0000000011111101",
								"0000000011010100",
								"0000000010100010",
								"0000000001111011",
								"0000000001010011",
								"0000000000110110",
								"0000000000001110",
								"1111111111101101",
								"1111111111000100",
								"1111111110100111",
								"1111111101111101",
								"1111111101100111",
								"1111111101001010",
								"1111111100111010",
								"1111111100100101",
								"1111111100100010",
								"1111111100001110",
								"1111111100000100",
								"1111111011110101",
								"1111111011101100",
								"1111111011100010",
								"1111111011100100",
								"1111111011110101",
								"1111111100010101",
								"1111111100111110",
								"1111111101100010",
								"1111111110000011",
								"1111111110010000",
								"1111111110000011",
								"1111111101111010",
								"1111111101101001",
								"1111111101101000",
								"1111111101111110",
								"1111111110100100",
								"1111111111100010",
								"0000000000100011",
								"0000000001011110",
								"0000000010001111",
								"0000000010100100",
								"0000000010101110",
								"0000000010011100",
								"0000000010010000",
								"0000000010000000",
								"0000000010000000",
								"0000000010000010",
								"0000000010010100",
								"0000000010101111",
								"0000000011010010",
								"0000000011101111",
								"0000000100001010",
								"0000000100011011",
								"0000000100100010",
								"0000000100110001",
								"0000000101001101",
								"0000000101100011",
								"0000000110000101",
								"0000000110010111",
								"0000000110111001",
								"0000000111000100",
								"0000000111001000",
								"0000000110101101",
								"0000000101110010",
								"0000000100101010",
								"0000000011010011",
								"0000000001111100",
								"0000000000101111",
								"1111111111110001",
								"1111111111001010",
								"1111111110110100",
								"1111111110100111",
								"1111111110010101",
								"1111111110000111",
								"1111111101101101",
								"1111111101001001",
								"1111111100001101",
								"1111111011010011",
								"1111111010101011",
								"1111111010000110",
								"1111111001111001",
								"1111111001110101",
								"1111111001111011",
								"1111111010000100",
								"1111111001110110",
								"1111111001011101",
								"1111111001000111",
								"1111111000101111",
								"1111111000100011",
								"1111111000011011",
								"1111111000101101",
								"1111111001000101",
								"1111111001101010",
								"1111111010011001",
								"1111111011001100",
								"1111111100000011",
								"1111111100111111",
								"1111111110000011",
								"1111111111001110",
								"0000000000011011",
								"0000000001100110",
								"0000000010100111",
								"0000000011011010",
								"0000000011110111",
								"0000000011111111",
								"0000000100000001",
								"0000000011110101",
								"0000000011110011",
								"0000000011111011",
								"0000000011111110",
								"0000000100010000",
								"0000000100011000",
								"0000000100101000",
								"0000000100101100",
								"0000000100101111",
								"0000000100101101",
								"0000000100011101",
								"0000000100010000",
								"0000000011111100",
								"0000000011100100",
								"0000000011001010",
								"0000000010110001",
								"0000000010101000",
								"0000000010101101",
								"0000000010111101",
								"0000000011011010",
								"0000000011111000",
								"0000000100001001",
								"0000000100001000",
								"0000000011110001",
								"0000000011000100",
								"0000000010010010",
								"0000000001100000",
								"0000000000110111",
								"0000000000010000",
								"1111111111111000",
								"1111111111011010",
								"1111111111000100",
								"1111111110100011",
								"1111111110000100",
								"1111111101101110",
								"1111111101001101",
								"1111111100111011",
								"1111111100011011",
								"1111111100010101",
								"1111111100000010",
								"1111111011111110",
								"1111111100000111",
								"1111111100001101",
								"1111111100100000",
								"1111111100101110",
								"1111111100111111",
								"1111111101001010",
								"1111111101001101",
								"1111111101000100",
								"1111111100110110",
								"1111111100111010",
								"1111111100110000",
								"1111111100000011",
								"1111111011111011",
								"1111111100000110",
								"1111111100001101",
								"1111111100100100",
								"1111111100111100",
								"1111111101101011",
								"1111111110011010",
								"1111111111001011",
								"1111111111100111",
								"0000000000000111",
								"0000000000010011",
								"0000000000011111",
								"0000000000100000",
								"0000000000001100",
								"1111111111111101",
								"1111111111100111",
								"1111111111010101",
								"1111111111001111",
								"1111111111010110",
								"1111111111101111",
								"0000000000011010",
								"0000000001010111",
								"0000000010001000",
								"0000000010110101",
								"0000000011010101",
								"0000000011100110",
								"0000000011100010",
								"0000000011100111",
								"0000000011011011",
								"0000000011011110",
								"0000000011101001",
								"0000000011110111",
								"0000000100000011",
								"0000000100001110",
								"0000000100010000",
								"0000000100000111",
								"0000000011111111",
								"0000000011101111",
								"0000000011101001",
								"0000000011100111",
								"0000000011100101",
								"0000000011101011",
								"0000000011111001",
								"0000000011111111",
								"0000000100001001",
								"0000000011111100",
								"0000000011110001",
								"0000000011011101",
								"0000000010111000",
								"0000000010001101",
								"0000000001011100",
								"0000000000011100",
								"1111111111101000",
								"1111111110111100",
								"1111111110010010",
								"1111111101110010",
								"1111111101000000",
								"1111111100011111",
								"1111111011110010",
								"1111111011001011",
								"1111111010011111",
								"1111111001111110",
								"1111111001100001",
								"1111111000111101",
								"1111111000011010",
								"1111110111110000",
								"1111110111001110",
								"1111110110110001",
								"1111110110110111",
								"1111110111011010",
								"1111111000011100",
								"1111111001011111",
								"1111111010100011",
								"1111111011011100",
								"1111111011111101",
								"1111111100010010",
								"1111111100100100",
								"1111111100100110",
								"1111111100101111",
								"1111111100110100",
								"1111111101011001",
								"1111111101111101",
								"1111111110110111",
								"1111111111111000",
								"0000000000111110",
								"0000000001110101",
								"0000000010011111",
								"0000000010110100",
								"0000000010111000",
								"0000000010110111",
								"0000000010101011",
								"0000000010111101",
								"0000000011011010",
								"0000000100010001",
								"0000000101010110",
								"0000000110010000",
								"0000000111010010",
								"0000001000000010",
								"0000001000100001",
								"0000001000110110",
								"0000001000101101",
								"0000001000101000",
								"0000001000010000",
								"0000000111111001",
								"0000000111010111",
								"0000000110110110",
								"0000000110001111",
								"0000000101100111",
								"0000000100111100",
								"0000000100010001",
								"0000000011011001",
								"0000000010101100",
								"0000000010001011",
								"0000000001101100",
								"0000000001011101",
								"0000000001000111",
								"0000000000110011",
								"0000000000010001",
								"1111111111101110",
								"1111111111000000",
								"1111111110010101",
								"1111111101101010",
								"1111111101001000",
								"1111111100110001",
								"1111111100011101",
								"1111111100010011",
								"1111111100001001",
								"1111111011110111",
								"1111111011101000",
								"1111111011001110",
								"1111111011000011",
								"1111111010110001",
								"1111111010110001",
								"1111111010111010",
								"1111111011001011",
								"1111111011100110",
								"1111111011111000",
								"1111111100010011",
								"1111111100110100",
								"1111111101101101",
								"1111111110011100",
								"1111111111011111",
								"0000000000001001",
								"0000000000110100",
								"0000000000111110",
								"0000000001000110",
								"0000000000101110",
								"0000000000010110",
								"1111111111111101",
								"1111111111111001",
								"0000000000001100",
								"0000000000100100",
								"0000000001001011",
								"0000000001011010",
								"0000000001101110",
								"0000000001100101",
								"0000000001011010",
								"0000000001000001",
								"0000000000101000",
								"0000000000011100",
								"0000000000100001",
								"0000000000101011",
								"0000000001000111",
								"0000000001011101",
								"0000000001110000",
								"0000000001111001",
								"0000000001110001",
								"0000000001001111",
								"0000000000100111",
								"1111111111111000",
								"1111111111001110",
								"1111111110111011",
								"1111111110110011",
								"1111111111000101",
								"1111111111001011",
								"1111111111010010",
								"1111111111001111",
								"1111111110111111",
								"1111111110101111",
								"1111111110101000",
								"1111111110101010",
								"1111111111001100",
								"1111111111111000",
								"0000000000110101",
								"0000000001101100",
								"0000000010001110",
								"0000000010101100",
								"0000000010100010",
								"0000000010000100",
								"0000000001010100",
								"0000000000001111",
								"1111111111001001",
								"1111111110001100",
								"1111111101101001",
								"1111111101100111",
								"1111111101110101",
								"1111111110010110",
								"1111111110110100",
								"1111111111000011",
								"1111111111000101",
								"1111111110110011",
								"1111111110011111",
								"1111111110001010",
								"1111111110000010",
								"1111111110001011",
								"1111111110100000",
								"1111111110110000",
								"1111111110110111",
								"1111111110101010",
								"1111111110010110",
								"1111111110001100",
								"1111111110001110",
								"1111111110011100",
								"1111111111000000",
								"1111111111110000",
								"0000000000011000",
								"0000000001000100",
								"0000000001001010",
								"0000000001010001",
								"0000000000100111",
								"0000000000001100",
								"1111111111011101",
								"1111111110111111",
								"1111111110111010",
								"1111111111000011",
								"1111111111101000",
								"0000000000011100",
								"0000000001000101",
								"0000000001101110",
								"0000000001111001",
								"0000000001111001",
								"0000000001101011",
								"0000000001011110",
								"0000000001010000",
								"0000000001010001",
								"0000000001100000",
								"0000000001111010",
								"0000000010100100",
								"0000000011001110",
								"0000000011111010",
								"0000000100010100",
								"0000000100100011",
								"0000000100100000",
								"0000000100010010",
								"0000000100000011",
								"0000000011100010",
								"0000000011011001",
								"0000000011010011",
								"0000000011011101",
								"0000000011110101",
								"0000000100001010",
								"0000000100011011",
								"0000000100100000",
								"0000000100001110",
								"0000000011101000",
								"0000000010111001",
								"0000000001111010",
								"0000000000111111",
								"0000000000000001",
								"1111111111010000",
								"1111111110100011",
								"1111111101110111",
								"1111111101001111",
								"1111111100101010",
								"1111111100001001",
								"1111111011111010",
								"1111111011110000",
								"1111111011110010",
								"1111111011111101",
								"1111111100000110",
								"1111111100010110",
								"1111111100011010",
								"1111111100011000",
								"1111111100001101",
								"1111111011111001",
								"1111111011100111",
								"1111111011010110",
								"1111111011010100",
								"1111111011010010",
								"1111111011010100",
								"1111111011011010",
								"1111111011011010",
								"1111111011010110",
								"1111111011010110",
								"1111111011000111",
								"1111111011001111",
								"1111111011010010",
								"1111111011100111",
								"1111111100001000",
								"1111111100111011",
								"1111111101111001",
								"1111111111000010",
								"0000000000000101",
								"0000000001000100",
								"0000000001100100",
								"0000000001101111",
								"0000000001011100",
								"0000000000111011",
								"0000000000001101",
								"1111111111100011",
								"1111111111000110",
								"1111111110111001",
								"1111111111010001",
								"1111111111111011",
								"0000000000110011",
								"0000000001110001",
								"0000000010011101",
								"0000000011001111",
								"0000000011100110",
								"0000000011110001",
								"0000000011110000",
								"0000000011011101",
								"0000000011001111",
								"0000000011000000",
								"0000000011000010",
								"0000000011000001",
								"0000000011010010",
								"0000000011100011",
								"0000000011111010",
								"0000000100000000",
								"0000000011111010",
								"0000000011100111",
								"0000000011000011",
								"0000000010011010",
								"0000000001011101",
								"0000000000101011",
								"1111111111100100",
								"1111111110110010",
								"1111111110001101",
								"1111111101111110",
								"1111111110000100",
								"1111111110010110",
								"1111111110101100",
								"1111111111000101",
								"1111111111010010",
								"1111111111010110",
								"1111111111010011",
								"1111111111001110",
								"1111111111001001",
								"1111111111001110",
								"1111111111010111",
								"1111111111100101",
								"1111111111110010",
								"1111111111111010",
								"1111111111101111",
								"1111111111011011",
								"1111111110111101",
								"1111111110010011",
								"1111111101110101",
								"1111111101000111",
								"1111111100111001",
								"1111111100101000",
								"1111111100111000",
								"1111111101000010",
								"1111111101011101",
								"1111111101101001",
								"1111111101110100",
								"1111111101110010",
								"1111111101110110",
								"1111111101111100",
								"1111111110001001",
								"1111111110100010",
								"1111111111001110",
								"1111111111111000",
								"0000000000010101",
								"0000000000100011",
								"0000000000010111",
								"0000000000001010",
								"1111111111110100",
								"1111111111110000",
								"1111111111110001",
								"0000000000001101",
								"0000000000101111",
								"0000000001100010",
								"0000000010001101",
								"0000000010101001",
								"0000000010101110",
								"0000000010010101",
								"0000000001111010",
								"0000000001010100",
								"0000000000110111",
								"0000000000101010",
								"0000000000100111",
								"0000000000110001",
								"0000000001000010",
								"0000000001001001",
								"0000000001010111",
								"0000000001010000",
								"0000000001001011",
								"0000000000101101",
								"0000000000010111",
								"1111111111101101",
								"1111111111001100",
								"1111111110100011",
								"1111111110001010",
								"1111111101110110",
								"1111111101101001",
								"1111111101011011",
								"1111111101001110",
								"1111111101000100",
								"1111111100111001",
								"1111111100111001",
								"1111111101000000",
								"1111111101010001",
								"1111111101101110",
								"1111111110100010",
								"1111111111010110",
								"0000000000000011",
								"0000000000100001",
								"0000000000101010",
								"0000000000011110",
								"0000000000001001",
								"1111111111100101",
								"1111111110111010",
								"1111111110100010",
								"1111111110010001",
								"1111111110100000",
								"1111111111001100",
								"0000000000000001",
								"0000000001010000",
								"0000000010001100",
								"0000000011001100",
								"0000000011101000",
								"0000000011110001",
								"0000000011011101",
								"0000000010111100",
								"0000000010100110",
								"0000000010010010",
								"0000000010010111",
								"0000000010011101",
								"0000000010111110",
								"0000000011001110",
								"0000000011101100",
								"0000000011110100",
								"0000000011111101",
								"0000000011011111",
								"0000000010101111",
								"0000000001011101",
								"1111111111111101",
								"1111111110101011",
								"1111111101101110",
								"1111111101100011",
								"1111111101111000",
								"1111111110101001",
								"1111111111110010",
								"0000000000011011",
								"0000000000110010",
								"0000000000010101",
								"1111111111100011",
								"1111111110001101",
								"1111111101000011",
								"1111111100001001",
								"1111111011011001",
								"1111111011001100",
								"1111111011001100",
								"1111111011101000",
								"1111111100000000",
								"1111111100011010",
								"1111111100100011",
								"1111111100101010",
								"1111111100100111",
								"1111111100100010",
								"1111111100101010",
								"1111111100101111",
								"1111111101000001",
								"1111111101011111",
								"1111111101110010",
								"1111111110010010",
								"1111111110101011",
								"1111111111000011",
								"1111111111011110",
								"1111111111110011",
								"0000000000011001",
								"0000000000110010",
								"0000000001011010",
								"0000000010000101",
								"0000000010101010",
								"0000000011001010",
								"0000000011010101",
								"0000000011010011",
								"0000000010111101",
								"0000000010100101",
								"0000000010000001",
								"0000000001101100",
								"0000000001100100",
								"0000000001100101",
								"0000000001110110",
								"0000000010001010",
								"0000000010101001",
								"0000000010110001",
								"0000000010110000",
								"0000000010010001",
								"0000000001100100",
								"0000000000101111",
								"1111111111111110",
								"1111111111011100",
								"1111111111001110",
								"1111111111001011",
								"1111111111010011",
								"1111111111011001",
								"1111111111011000",
								"1111111111000111",
								"1111111110100000",
								"1111111101101000",
								"1111111100101010",
								"1111111011110101",
								"1111111011010100",
								"1111111011001010",
								"1111111011100011",
								"1111111100001010",
								"1111111101000001",
								"1111111110000011",
								"1111111110110111",
								"1111111111100110",
								"0000000000000000",
								"0000000000001001",
								"0000000000001000",
								"1111111111111011",
								"1111111111100111",
								"1111111111010011",
								"1111111111000110",
								"1111111111000110",
								"1111111111011001",
								"1111111111110100",
								"0000000000100010",
								"0000000001000011",
								"0000000001100110",
								"0000000010000000",
								"0000000010010011",
								"0000000010011011",
								"0000000010011011",
								"0000000010010011",
								"0000000010000101",
								"0000000010000100",
								"0000000010001000",
								"0000000010011111",
								"0000000011000000",
								"0000000011011111"
								);
								
	variable expected_out : WAV_IN := ("0000000011001100",
									"0000000110110100",
									"0000001001110100",
									"0000001100111011",
									"0000001100100011",
									"0000001100001001",
									"0000001100011110",
									"0000001101010110",
									"0000001110110100",
									"0000010000011101",
									"0000010001111010",
									"0000010010110011",
									"0000010010111001",
									"0000010001110111",
									"0000010000000111",
									"0000001101101001",
									"0000001010111111",
									"0000001000011110",
									"0000000110011100",
									"0000000101000001",
									"0000000100001100",
									"0000000011110110",
									"0000000011101111",
									"0000000011101000",
									"0000000011010010",
									"0000000010011100",
									"0000000001001000",
									"1111111111010001",
									"1111111101000110",
									"1111111010110011",
									"1111111000101100",
									"1111110110110101",
									"1111110101011111",
									"1111110100101100",
									"1111110100010101",
									"1111110100100101",
									"1111110101010000",
									"1111110110010010",
									"1111110111100100",
									"1111111000100011",
									"1111111001010110",
									"1111111001100001",
									"1111111001011001",
									"1111111001000100",
									"1111111000101100",
									"1111111000101101",
									"1111111000111010",
									"1111111001100110",
									"1111111010011110",
									"1111111011010101",
									"1111111011111010",
									"1111111100000000",
									"1111111011011110",
									"1111111010010001",
									"1111111000110000",
									"1111110111000101",
									"1111110101101110",
									"1111110101000001",
									"1111110100110101",
									"1111110101100110",
									"1111110110111011",
									"1111111000111101",
									"1111111011011011",
									"1111111110000010",
									"0000000000100110",
									"0000000010100110",
									"0000000100000000",
									"0000000100011100",
									"0000000100000010",
									"0000000010111110",
									"0000000001100001",
									"1111111111110001",
									"1111111110001110",
									"1111111100111101",
									"1111111100010101",
									"1111111100101001",
									"1111111101100111",
									"1111111111010100",
									"0000000001001110",
									"0000000011000001",
									"0000000100100110",
									"0000000101100101",
									"0000000110001101",
									"0000000110100010",
									"0000000110100111",
									"0000000110101101",
									"0000000110100101",
									"0000000110010101",
									"0000000101110100",
									"0000000101000110",
									"0000000100001001",
									"0000000011001001",
									"0000000010010001",
									"0000000001100011",
									"0000000001010100",
									"0000000001010111",
									"0000000001110001",
									"0000000010010001",
									"0000000010101011",
									"0000000010111111",
									"0000000010111000",
									"0000000010100100",
									"0000000001111011",
									"0000000001001110",
									"0000000000101110",
									"0000000000100100",
									"0000000001000000",
									"0000000001110110",
									"0000000011000110",
									"0000000100010110",
									"0000000101100110",
									"0000000110100001",
									"0000000111001001",
									"0000000111100011",
									"0000000111101101",
									"0000000111100110",
									"0000000111001100",
									"0000000110011111",
									"0000000101100010",
									"0000000100101000",
									"0000000011101110",
									"0000000011001101",
									"0000000010111010",
									"0000000011000111",
									"0000000011101011",
									"0000000100100000",
									"0000000101011000",
									"0000000110000011",
									"0000000110011110",
									"0000000110100100",
									"0000000110011001",
									"0000000110010001",
									"0000000110001010",
									"0000000101111110",
									"0000000101110110",
									"0000000101010101",
									"0000000100101111",
									"0000000100000010",
									"0000000011101011",
									"0000000011101010",
									"0000000100001101",
									"0000000101001000",
									"0000000110001010",
									"0000000111000111",
									"0000000111100101",
									"0000000111100100",
									"0000000110111100",
									"0000000110000011",
									"0000000100111111",
									"0000000100001010",
									"0000000011100010",
									"0000000011000000",
									"0000000010100010",
									"0000000001110000",
									"0000000000100101",
									"1111111111000010",
									"1111111101001101",
									"1111111011010010",
									"1111111001101000",
									"1111111000001101",
									"1111110111000000",
									"1111110110011001",
									"1111110110001010",
									"1111110110100010",
									"1111110111001010",
									"1111110111110010",
									"1111110111111100",
									"1111110111100011",
									"1111110110101111",
									"1111110101011111",
									"1111110100010011",
									"1111110011010100",
									"1111110010110011",
									"1111110010110111",
									"1111110011101110",
									"1111110101010101",
									"1111110111110011",
									"1111111010110100",
									"1111111101111110",
									"0000000000110100",
									"0000000010111101",
									"0000000011111100",
									"0000000011111111",
									"0000000011000010",
									"0000000001011000",
									"1111111111101001",
									"1111111101111001",
									"1111111100100110",
									"1111111011110000",
									"1111111011010010",
									"1111111010111101",
									"1111111010110000",
									"1111111010101100",
									"1111111010110011",
									"1111111011011110",
									"1111111100100101",
									"1111111110000000",
									"1111111111101011",
									"0000000001011011",
									"0000000011001000",
									"0000000100100101",
									"0000000101011111",
									"0000000101011011",
									"0000000100011000",
									"0000000010101111",
									"0000000001001110",
									"0000000000010001",
									"0000000000001011",
									"0000000000110110",
									"0000000010001011",
									"0000000100001000",
									"0000000110101010",
									"0000001001110100",
									"0000001101000111",
									"0000010000011111",
									"0000010011001100",
									"0000010100100011",
									"0000010100011101",
									"0000010010010110",
									"0000001111010010",
									"0000001011100111",
									"0000001000011111",
									"0000000110011101",
									"0000000101100110",
									"0000000110000110",
									"0000000110111011",
									"0000000111110000",
									"0000000111100101",
									"0000000110000111",
									"0000000011111000",
									"0000000001001101",
									"1111111111000111",
									"1111111110001001",
									"1111111101101101",
									"1111111110001011",
									"1111111110101011",
									"1111111111001000",
									"1111111111100100",
									"1111111111011101",
									"1111111111011001",
									"1111111110110101",
									"1111111110001101",
									"1111111101100110",
									"1111111100111011",
									"1111111100101001",
									"1111111100100000",
									"1111111100101001",
									"1111111100111001",
									"1111111101001100",
									"1111111101100000",
									"1111111101111000",
									"1111111110010100",
									"1111111110110010",
									"1111111111011000",
									"0000000000000001",
									"0000000000111000",
									"0000000001110010",
									"0000000010110111",
									"0000000011101010",
									"0000000100000110",
									"0000000011111000",
									"0000000011000001",
									"0000000001101110",
									"0000000000010110",
									"1111111111100010",
									"1111111111010011",
									"0000000000000110",
									"0000000001011110",
									"0000000011000000",
									"0000000100100000",
									"0000000101010001",
									"0000000101001101",
									"0000000100011100",
									"0000000011000100",
									"0000000001101101",
									"0000000000101110",
									"0000000000011001",
									"0000000000111010",
									"0000000010010011",
									"0000000100011000",
									"0000000111000111",
									"0000001010000110",
									"0000001100101101",
									"0000001110101010",
									"0000001111001111",
									"0000001110011000",
									"0000001100001001",
									"0000001000110000",
									"0000000101000010",
									"0000000001011101",
									"1111111110011111",
									"1111111100011111",
									"1111111011010000",
									"1111111010011101",
									"1111111001111010",
									"1111111001000110",
									"1111110111111111",
									"1111110110100000",
									"1111110100101101",
									"1111110010111110",
									"1111110001001000",
									"1111101111100100",
									"1111101110011001",
									"1111101101100111",
									"1111101101100011",
									"1111101110001101",
									"1111101111101001",
									"1111110001110001",
									"1111110100010010",
									"1111110110111100",
									"1111111001011010",
									"1111111011101110",
									"1111111101111100",
									"0000000000001011",
									"0000000010011010",
									"0000000100101011",
									"0000000110110001",
									"0000001000101011",
									"0000001010011000",
									"0000001011110000",
									"0000001100110101",
									"0000001101110001",
									"0000001110100111",
									"0000001111010111",
									"0000010000001101",
									"0000010000111001",
									"0000010001011001",
									"0000010001011001",
									"0000010000110000",
									"0000001111010100",
									"0000001101010110",
									"0000001011001000",
									"0000001001001101",
									"0000001000001000",
									"0000000111110000",
									"0000001000001010",
									"0000001000110010",
									"0000001000110111",
									"0000001000001101",
									"0000000110010100",
									"0000000011011001",
									"1111111111111001",
									"1111111100001110",
									"1111111001001100",
									"1111110111000001",
									"1111110110000011",
									"1111110110000010",
									"1111110110100110",
									"1111110111010100",
									"1111110111101110",
									"1111110111101010",
									"1111110110111011",
									"1111110101101001",
									"1111110011111100",
									"1111110010000110",
									"1111110000011010",
									"1111101111001010",
									"1111101110001000",
									"1111101101000101",
									"1111101011111101",
									"1111101010011010",
									"1111101000110100",
									"1111100111001000",
									"1111100101100111",
									"1111100100100100",
									"1111100100001110",
									"1111100101010101",
									"1111100111101111",
									"1111101011100100",
									"1111110000010101",
									"1111110101011000",
									"1111111010010001",
									"1111111110011010",
									"0000000001100010",
									"0000000011101010",
									"0000000101000110",
									"0000000110001001",
									"0000000111010000",
									"0000001000101110",
									"0000001010110110",
									"0000001101101010",
									"0000010000101100",
									"0000010011101111",
									"0000010110000011",
									"0000010111100001",
									"0000011000010001",
									"0000011000010011",
									"0000011000010110",
									"0000011000101110",
									"0000011001100010",
									"0000011010110111",
									"0000011100001010",
									"0000011101001100",
									"0000011101100110",
									"0000011101010000",
									"0000011100001001",
									"0000011010001011",
									"0000010111101100",
									"0000010100101110",
									"0000010001011001",
									"0000001101101111",
									"0000001001101101",
									"0000000101010101",
									"0000000000101110",
									"1111111100001010",
									"1111110111111110",
									"1111110100100010",
									"1111110010001001",
									"1111110000101111",
									"1111110000010100",
									"1111110000011000",
									"1111110000011100",
									"1111110000011111",
									"1111110000000100",
									"1111101111011111",
									"1111101110110010",
									"1111101110000100",
									"1111101101100101",
									"1111101101010000",
									"1111101101011011",
									"1111101101110111",
									"1111101110101010",
									"1111101111110011",
									"1111110001000110",
									"1111110010100101",
									"1111110011111001",
									"1111110100110000",
									"1111110100111101",
									"1111110100010100",
									"1111110011000100",
									"1111110001101000",
									"1111110000011101",
									"1111110000000110",
									"1111110000111010",
									"1111110010110001",
									"1111110101011001",
									"1111111000010011",
									"1111111011000111",
									"1111111101100001",
									"1111111111100111",
									"0000000001011010",
									"0000000011000111",
									"0000000100111011",
									"0000000110100111",
									"0000001000011110",
									"0000001010000110",
									"0000001011101111",
									"0000001101001000",
									"0000001110010011",
									"0000001111010000",
									"0000001111100100",
									"0000001111101100",
									"0000001111001110",
									"0000001110011110",
									"0000001101100110",
									"0000001100101001",
									"0000001011111100",
									"0000001011100110",
									"0000001011101111",
									"0000001011111111",
									"0000001100011100",
									"0000001101011101",
									"0000001110011000",
									"0000001111001100",
									"0000001111101111",
									"0000001111001110",
									"0000001110001101",
									"0000001100101000",
									"0000001010011011",
									"0000000111110100",
									"0000000101001001",
									"0000000010101101",
									"0000000000110100",
									"1111111111100000",
									"1111111110100111",
									"1111111110100010",
									"1111111110111000",
									"1111111111110000",
									"0000000000111011",
									"0000000001111000",
									"0000000010011111",
									"0000000010010111",
									"0000000001010010",
									"1111111111001010",
									"1111111100011000",
									"1111111001010010",
									"1111110110010111",
									"1111110100001000",
									"1111110010101110",
									"1111110001111100",
									"1111110001110110",
									"1111110001111110",
									"1111110001110111",
									"1111110001100111",
									"1111110000111111",
									"1111110000001111",
									"1111101111101000",
									"1111101111011000",
									"1111101111011100",
									"1111101111111011",
									"1111110000100010",
									"1111110001000010",
									"1111110001011100",
									"1111110001100000",
									"1111110001010000",
									"1111110000111000",
									"1111110000010100",
									"1111110000000011",
									"1111110000001011",
									"1111110000101101",
									"1111110001111110",
									"1111110011101101",
									"1111110110000010",
									"1111111001000011",
									"1111111100010011",
									"1111111111100100",
									"0000000010101110",
									"0000000101011000",
									"0000001000000000",
									"0000001010011101",
									"0000001100111101",
									"0000001111100100",
									"0000010010000101",
									"0000010100100110",
									"0000010110110111",
									"0000011001000101",
									"0000011011001010",
									"0000011101011000",
									"0000011111101011",
									"0000100001110111",
									"0000100011011010",
									"0000100011110000",
									"0000100010100010",
									"0000011111110100",
									"0000011100001000",
									"0000011000000110",
									"0000010100100101",
									"0000010001110010",
									"0000001111110001",
									"0000001110100111",
									"0000001101110101",
									"0000001101010011",
									"0000001100011110",
									"0000001011000111",
									"0000001000111111",
									"0000000101111011",
									"0000000010010110",
									"1111111110011110",
									"1111111010110110",
									"1111110111111010",
									"1111110110000000",
									"1111110100111110",
									"1111110100110010",
									"1111110100101001",
									"1111110100000111",
									"1111110010101101",
									"1111110000000010",
									"1111101100101111",
									"1111101000110111",
									"1111100101000110",
									"1111100001111011",
									"1111011111010101",
									"1111011101111010",
									"1111011101010100",
									"1111011101100101",
									"1111011110100010",
									"1111011111111000",
									"1111100001101010",
									"1111100011101011",
									"1111100101111101",
									"1111101000011000",
									"1111101010111101",
									"1111101101110011",
									"1111110000101110",
									"1111110011011111",
									"1111110110000100",
									"1111111000000000",
									"1111111001100101",
									"1111111010111101",
									"1111111100011000",
									"1111111110000111",
									"0000000000001110",
									"0000000010101100",
									"0000000101010011",
									"0000000111111001",
									"0000001010001000",
									"0000001100000000",
									"0000001101010111",
									"0000001110010110",
									"0000001111010000",
									"0000010000000101",
									"0000010001001010",
									"0000010010010000",
									"0000010011010110",
									"0000010100001101",
									"0000010100100001",
									"0000010100011001",
									"0000010011100100",
									"0000010010011101",
									"0000010001000100",
									"0000001111011011",
									"0000001101010100",
									"0000001010110000",
									"0000000111100100",
									"0000000100001111",
									"0000000001001000",
									"1111111110100110",
									"1111111100111111",
									"1111111100011010",
									"1111111100111000",
									"1111111101111001",
									"1111111111000110",
									"1111111111101000",
									"1111111111011010",
									"1111111110001100",
									"1111111100101011",
									"1111111011001001",
									"1111111010001000",
									"1111111001111001",
									"1111111010010010",
									"1111111011011000",
									"1111111100100001",
									"1111111101011010",
									"1111111101110000",
									"1111111101010001",
									"1111111100010000",
									"1111111011000001",
									"1111111001110011",
									"1111111001001001",
									"1111111001010111",
									"1111111010100000",
									"1111111100100001",
									"1111111111000100",
									"0000000001011000",
									"0000000011001100",
									"0000000011111111",
									"0000000100000010",
									"0000000011101011",
									"0000000011001111",
									"0000000011010101",
									"0000000011110001",
									"0000000100011011",
									"0000000101000000",
									"0000000100110011",
									"0000000011101010",
									"0000000001011101",
									"1111111110011011",
									"1111111011011001",
									"1111111000100101",
									"1111110110111000",
									"1111110110100000",
									"1111110111011010",
									"1111111001110111",
									"1111111101010000",
									"0000000001001000",
									"0000000100110011",
									"0000000111011011",
									"0000001000101111",
									"0000001000100101",
									"0000000111011010",
									"0000000101111110",
									"0000000100101110",
									"0000000100010001",
									"0000000100100110",
									"0000000101011111",
									"0000000110100010",
									"0000000111001010",
									"0000000111001001",
									"0000000110100011",
									"0000000101101110",
									"0000000101001111",
									"0000000101011001",
									"0000000101111101",
									"0000000110100110",
									"0000000110110100",
									"0000000110001010",
									"0000000100100110",
									"0000000010011100",
									"1111111111110100",
									"1111111101101010",
									"1111111100001001",
									"1111111011111010",
									"1111111100110010",
									"1111111110011111",
									"0000000000110001",
									"0000000010011110",
									"0000000011100111",
									"0000000011011100",
									"0000000001111111",
									"1111111111110100",
									"1111111101001001",
									"1111111010111000",
									"1111111001011011",
									"1111111000110101",
									"1111111001000101",
									"1111111001101110",
									"1111111010010110",
									"1111111010100001",
									"1111111010000101",
									"1111111000110001",
									"1111110110110100",
									"1111110100011010",
									"1111110010000000",
									"1111110000000001",
									"1111101110101111",
									"1111101110010111",
									"1111101110101000",
									"1111101111101001",
									"1111110000110000",
									"1111110001101111",
									"1111110010010101",
									"1111110010000010",
									"1111110001010001",
									"1111110000001001",
									"1111101111000110",
									"1111101110101101",
									"1111101111001111",
									"1111110000110001",
									"1111110011010111",
									"1111110110100110",
									"1111111010001101",
									"1111111101110110",
									"0000000001001101",
									"0000000100010101",
									"0000000111000111",
									"0000001001101101",
									"0000001100000111",
									"0000001110000100",
									"0000001111100011",
									"0000010000011011",
									"0000010000100111",
									"0000010000011011",
									"0000001111110101",
									"0000001111001101",
									"0000001110110010",
									"0000001110101011",
									"0000001111001000",
									"0000001111111011",
									"0000010000111101",
									"0000010001110110",
									"0000010010011101",
									"0000010010110000",
									"0000010010101100",
									"0000010010100110",
									"0000010010100010",
									"0000010010100000",
									"0000010010110011",
									"0000010010111110",
									"0000010011000010",
									"0000010010110001",
									"0000010001110000",
									"0000010000000100",
									"0000001101011101",
									"0000001010000010",
									"0000000110000101",
									"0000000001111100",
									"1111111110010001",
									"1111111011100100",
									"1111111010001101",
									"1111111010010110",
									"1111111011101101",
									"1111111101111001",
									"0000000000001111",
									"0000000010010001",
									"0000000011001101",
									"0000000010110101",
									"0000000001001000",
									"1111111110010000",
									"1111111011000100",
									"1111110111110000",
									"1111110100111101",
									"1111110010111101",
									"1111110001101010",
									"1111110001011100",
									"1111110001110011",
									"1111110010100100",
									"1111110011010010",
									"1111110011101110",
									"1111110011101011",
									"1111110011001000",
									"1111110010010000",
									"1111110001010001",
									"1111110000101001",
									"1111110000100101",
									"1111110001011100",
									"1111110011000010",
									"1111110101011111",
									"1111111000011011",
									"1111111011111010",
									"1111111111100010",
									"0000000010110010",
									"0000000101011111",
									"0000000110111111",
									"0000000111011011",
									"0000000110111100",
									"0000000101110101",
									"0000000100100111",
									"0000000011100111",
									"0000000011000000",
									"0000000010110111",
									"0000000011000000",
									"0000000011001000",
									"0000000011000100",
									"0000000010101101",
									"0000000010000100",
									"0000000001011000",
									"0000000001000000",
									"0000000001001010",
									"0000000001111111",
									"0000000011100110",
									"0000000101100000",
									"0000000111110100",
									"0000001001111000",
									"0000001011100011",
									"0000001100100000",
									"0000001100100101",
									"0000001100000001",
									"0000001011000000",
									"0000001010000100",
									"0000001001010100",
									"0000001000111011",
									"0000001000101000",
									"0000001000010011",
									"0000000111100011",
									"0000000110001011",
									"0000000100001111",
									"0000000010000011",
									"0000000000000010",
									"1111111110111001",
									"1111111110100111",
									"1111111111001000",
									"1111111111111011",
									"0000000000100001",
									"0000000000011110",
									"1111111111100011",
									"1111111101110001",
									"1111111011010101",
									"1111111000111001",
									"1111110110111010",
									"1111110110000111",
									"1111110110011010",
									"1111110111101111",
									"1111111001100110",
									"1111111011010001",
									"1111111100100100",
									"1111111101000111",
									"1111111100111100",
									"1111111100011101",
									"1111111011101101",
									"1111111011001110",
									"1111111011000101",
									"1111111011100001",
									"1111111100100001",
									"1111111110000100",
									"0000000000000011",
									"0000000010001101",
									"0000000100011010",
									"0000000110010001",
									"0000000111110100",
									"0000001000111100",
									"0000001001111000",
									"0000001010101010",
									"0000001011011010",
									"0000001011111100",
									"0000001100001010",
									"0000001011111101",
									"0000001011001000",
									"0000001001011111",
									"0000000111001001",
									"0000000100010111",
									"0000000001100100",
									"1111111111011100",
									"1111111110010100",
									"1111111110001110",
									"1111111111001010",
									"0000000000111010",
									"0000000010110110",
									"0000000100101110",
									"0000000101110011",
									"0000000101100001",
									"0000000100000010",
									"0000000001000011",
									"1111111101010111",
									"1111111001010111",
									"1111110101110000",
									"1111110011001111",
									"1111110001111110",
									"1111110010001110",
									"1111110011010000",
									"1111110100101111",
									"1111110101110101",
									"1111110110010100",
									"1111110101111100",
									"1111110101000000",
									"1111110011101011",
									"1111110010010100",
									"1111110001010101",
									"1111110001000100",
									"1111110010000001",
									"1111110100011000",
									"1111111000011000",
									"1111111101001100",
									"0000000010001101",
									"0000000110000111",
									"0000001000001100",
									"0000001000001110",
									"0000000110001010",
									"0000000011010010",
									"0000000000011000",
									"1111111110101100",
									"1111111110111011",
									"0000000001001001",
									"0000000100111000",
									"0000001001000100",
									"0000001101001110",
									"0000010000001111",
									"0000010010000110",
									"0000010010100111",
									"0000010010000000",
									"0000010000110010",
									"0000001111011011",
									"0000001110011001",
									"0000001101110010",
									"0000001101101010",
									"0000001101100011",
									"0000001101011110",
									"0000001101000100",
									"0000001100000111",
									"0000001010111111",
									"0000001001011100",
									"0000000111110010",
									"0000000110001110",
									"0000000100100010",
									"0000000011000001",
									"0000000001010011",
									"1111111111100100",
									"1111111101101000",
									"1111111011010110",
									"1111111001000101",
									"1111110110101101",
									"1111110100110010",
									"1111110011100100",
									"1111110011010001",
									"1111110011110110",
									"1111110101001010",
									"1111110110110001",
									"1111111000001010",
									"1111111001001010",
									"1111111001010101",
									"1111111000110111",
									"1111110111110010",
									"1111110110100110",
									"1111110101101100",
									"1111110101100101",
									"1111110110101010",
									"1111111000101100",
									"1111111011011110",
									"1111111110010011",
									"0000000000101001",
									"0000000010001101",
									"0000000010111000",
									"0000000010111011",
									"0000000010110001",
									"0000000010110101",
									"0000000011101000",
									"0000000101011001",
									"0000001000000111",
									"0000001011011001",
									"0000001110100101",
									"0000010001000011",
									"0000010010001010",
									"0000010001110101",
									"0000010000001000",
									"0000001101001111",
									"0000001001111011",
									"0000000110011111",
									"0000000011100000",
									"0000000001011010",
									"0000000000001001",
									"1111111111110100",
									"0000000000001101",
									"0000000001000011",
									"0000000010000101",
									"0000000010111010",
									"0000000011001000",
									"0000000010100111",
									"0000000001001011",
									"1111111111001110",
									"1111111101000001",
									"1111111010110101",
									"1111111001000100",
									"1111110111101100",
									"1111110110110111",
									"1111110110100100",
									"1111110110110010",
									"1111110111001001",
									"1111110111011100",
									"1111110111010000",
									"1111110110010101",
									"1111110100111010"
									);
	
	
	begin
		
		rst_l <= '0';
		wait until clk'event and clk='1';
		rst_l <= '1'; 
		
		for i in 0 to SAMPLES-1 loop	
			
			sample <= input(i);
			expected <= expected_out(i);
			
			
			wait until clk'event and clk='1'; 

			assert (output = expected)
			report "Mismatch for index i = " & integer'image(i)
			severity error;
			
		end loop;	 
		
		enable <= '0';
		end process;

end TB_Arch;

